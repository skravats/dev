module const_signals(
	output wire high,
	output wire low
);

assign high = 1'b1;
assign low  = 1'b0;

endmodule