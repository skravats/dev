// system_bd.v

// Generated using ACDS version 18.1.2 277

`timescale 1 ps / 1 ps
module system_bd (
		input  wire        tx_ref_clk_clk,                 //                 tx_ref_clk.clk
		input  wire        rx_ref_clk_clk,                 //                 rx_ref_clk.clk
		input  wire        tx_fifo_bypass_bypass,          //             tx_fifo_bypass.bypass
		input  wire        sys_clk_clk,                    //                    sys_clk.clk
		input  wire        sys_rst_reset_n,                //                    sys_rst.reset_n
		input  wire        sys_ddr3_cntrl_pll_ref_clk_clk, // sys_ddr3_cntrl_pll_ref_clk.clk
		input  wire        sys_ddr3_cntrl_oct_oct_rzqin,   //         sys_ddr3_cntrl_oct.oct_rzqin
		output wire [0:0]  sys_ddr3_cntrl_mem_mem_ck,      //         sys_ddr3_cntrl_mem.mem_ck
		output wire [0:0]  sys_ddr3_cntrl_mem_mem_ck_n,    //                           .mem_ck_n
		output wire [11:0] sys_ddr3_cntrl_mem_mem_a,       //                           .mem_a
		output wire [2:0]  sys_ddr3_cntrl_mem_mem_ba,      //                           .mem_ba
		output wire [0:0]  sys_ddr3_cntrl_mem_mem_cke,     //                           .mem_cke
		output wire [0:0]  sys_ddr3_cntrl_mem_mem_cs_n,    //                           .mem_cs_n
		output wire [0:0]  sys_ddr3_cntrl_mem_mem_odt,     //                           .mem_odt
		output wire [0:0]  sys_ddr3_cntrl_mem_mem_reset_n, //                           .mem_reset_n
		output wire [0:0]  sys_ddr3_cntrl_mem_mem_we_n,    //                           .mem_we_n
		output wire [0:0]  sys_ddr3_cntrl_mem_mem_ras_n,   //                           .mem_ras_n
		output wire [0:0]  sys_ddr3_cntrl_mem_mem_cas_n,   //                           .mem_cas_n
		inout  wire [7:0]  sys_ddr3_cntrl_mem_mem_dqs,     //                           .mem_dqs
		inout  wire [7:0]  sys_ddr3_cntrl_mem_mem_dqs_n,   //                           .mem_dqs_n
		inout  wire [63:0] sys_ddr3_cntrl_mem_mem_dq,      //                           .mem_dq
		output wire [7:0]  sys_ddr3_cntrl_mem_mem_dm,      //                           .mem_dm
		output wire        sys_ethernet_mdio_mdc,          //          sys_ethernet_mdio.mdc
		input  wire        sys_ethernet_mdio_mdio_in,      //                           .mdio_in
		output wire        sys_ethernet_mdio_mdio_out,     //                           .mdio_out
		output wire        sys_ethernet_mdio_mdio_oen,     //                           .mdio_oen
		input  wire        sys_ethernet_ref_clk_clk,       //       sys_ethernet_ref_clk.clk
		input  wire        sys_ethernet_sgmii_rxp_0,       //         sys_ethernet_sgmii.rxp_0
		output wire        sys_ethernet_sgmii_txp_0,       //                           .txp_0
		output wire        sys_ethernet_reset_reset,       //         sys_ethernet_reset.reset
		output wire [23:0] sys_flash_tcm_address_out,      //                  sys_flash.tcm_address_out
		output wire [0:0]  sys_flash_tcm_read_n_out,       //                           .tcm_read_n_out
		output wire [0:0]  sys_flash_tcm_write_n_out,      //                           .tcm_write_n_out
		inout  wire [31:0] sys_flash_tcm_data_out,         //                           .tcm_data_out
		output wire [0:0]  sys_flash_tcm_chipselect_n_out, //                           .tcm_chipselect_n_out
		input  wire [31:0] sys_gpio_bd_in_port,            //                sys_gpio_bd.in_port
		output wire [31:0] sys_gpio_bd_out_port,           //                           .out_port
		input  wire [31:0] sys_gpio_in_export,             //                sys_gpio_in.export
		output wire [31:0] sys_gpio_out_export,            //               sys_gpio_out.export
		input  wire        sys_spi_MISO,                   //                    sys_spi.MISO
		output wire        sys_spi_MOSI,                   //                           .MOSI
		output wire        sys_spi_SCLK,                   //                           .SCLK
		output wire [7:0]  sys_spi_SS_n                    //                           .SS_n
	);

	wire          sys_clk_clk_clk;                                                    // sys_clk:clk_out -> [ad9144_jesd204:sys_clk_clk, ad9680_jesd204:sys_clk_clk, avalon_st_adapter:in_clk_0_clk, avalon_st_adapter_001:in_clk_0_clk, avl_adxcfg_0:rcfg_clk, avl_adxcfg_1:rcfg_clk, avl_adxcfg_2:rcfg_clk, avl_adxcfg_3:rcfg_clk, axi_ad9144_dma:s_axi_aclk, axi_ad9680_dma:s_axi_aclk, irq_mapper:clk, mm_interconnect_0:sys_clk_clk_clk, mm_interconnect_1:sys_clk_clk_clk, mm_interconnect_2:sys_clk_clk_clk, rst_controller:clk, rst_controller_004:clk, rst_controller_005:clk, sys_cpu:clk, sys_ethernet:clk, sys_ethernet:ff_rx_clk, sys_ethernet:ff_tx_clk, sys_ethernet_dma_rx:clock_clk, sys_ethernet_dma_tx:clock_clk, sys_ethernet_reset:clk, sys_flash:clk_clk, sys_flash_bridge:clk, sys_gpio_bd:clk, sys_gpio_in:clk, sys_gpio_out:clk, sys_id:clock, sys_int_mem:clk, sys_spi:clk, sys_timer_1:clk, sys_timer_2:clk, sys_tlb_mem:clk, sys_tlb_mem:clk2, sys_uart:clk]
	wire          sys_dma_clk_clk_clk;                                                // sys_dma_clk:clk_out -> [ad9680_adcfifo:dma_clk, avl_ad9144_fifo:dma_clk, axi_ad9144_dma:m_axis_aclk, axi_ad9144_dma:m_src_axi_aclk, axi_ad9680_dma:m_dest_axi_aclk, axi_ad9680_dma:s_axis_aclk]
	wire          sys_ddr3_cntrl_emif_usr_clk_clk;                                    // sys_ddr3_cntrl:emif_usr_clk -> [mm_interconnect_0:sys_ddr3_cntrl_emif_usr_clk_clk, rst_controller_002:clk, rst_controller_006:clk, sys_dma_clk:in_clk]
	wire          ad9680_jesd204_link_clk_clk;                                        // ad9680_jesd204:link_clk_clk -> [ad9680_adcfifo:adc_clk, rst_controller_001:clk]
	wire          ad9144_jesd204_link_clk_clk;                                        // ad9144_jesd204:link_clk_clk -> [avl_ad9144_fifo:dac_clk, rst_controller_003:clk, util_ad9144_upack:dac_clk]
	wire  [127:0] avl_ad9144_fifo_if_dac_data_data;                                   // avl_ad9144_fifo:dac_data -> util_ad9144_upack:dac_data
	wire          util_ad9144_upack_if_dac_valid_valid;                               // util_ad9144_upack:dac_valid -> avl_ad9144_fifo:dac_valid
	wire          avl_ad9144_fifo_if_dma_ready_ready;                                 // avl_ad9144_fifo:dma_ready -> axi_ad9144_dma:m_axis_ready
	wire  [127:0] ad9680_adcfifo_if_dma_wdata_data;                                   // ad9680_adcfifo:dma_wdata -> axi_ad9680_dma:s_axis_data
	wire          ad9680_adcfifo_if_dma_wr_valid;                                     // ad9680_adcfifo:dma_wr -> axi_ad9680_dma:s_axis_valid
	wire          axi_ad9680_dma_if_s_axis_ready_ready;                               // axi_ad9680_dma:s_axis_ready -> ad9680_adcfifo:dma_wready
	wire          axi_ad9680_dma_if_s_axis_xfer_req_xfer_req;                         // axi_ad9680_dma:s_axis_xfer_req -> ad9680_adcfifo:dma_xfer_req
	wire  [127:0] axi_ad9144_dma_if_m_axis_data_data;                                 // axi_ad9144_dma:m_axis_data -> avl_ad9144_fifo:dma_data
	wire          axi_ad9144_dma_if_m_axis_last_last;                                 // axi_ad9144_dma:m_axis_last -> avl_ad9144_fifo:dma_xfer_last
	wire          axi_ad9144_dma_if_m_axis_valid_valid;                               // axi_ad9144_dma:m_axis_valid -> avl_ad9144_fifo:dma_valid
	wire          axi_ad9144_dma_if_m_axis_xfer_req_xfer_req;                         // axi_ad9144_dma:m_axis_xfer_req -> avl_ad9144_fifo:dma_xfer_req
	wire          sys_clk_clk_reset_reset;                                            // sys_clk:reset_n_out -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_004:reset_in0, rst_controller_005:reset_in0, sys_ddr3_cntrl:global_reset_n]
	wire          sys_ddr3_cntrl_emif_usr_reset_n_reset;                              // sys_ddr3_cntrl:emif_usr_reset_n -> [rst_controller_006:reset_in0, sys_dma_clk:reset_n]
	wire          sys_flash_tcm_data_outen;                                           // sys_flash:tcm_data_outen -> sys_flash_bridge:tcs_tcm_data_outen
	wire          sys_flash_tcm_request;                                              // sys_flash:tcm_request -> sys_flash_bridge:request
	wire          sys_flash_tcm_write_n_out_signal;                                   // sys_flash:tcm_write_n_out -> sys_flash_bridge:tcs_tcm_write_n_out
	wire          sys_flash_tcm_read_n_out_signal;                                    // sys_flash:tcm_read_n_out -> sys_flash_bridge:tcs_tcm_read_n_out
	wire          sys_flash_tcm_grant;                                                // sys_flash_bridge:grant -> sys_flash:tcm_grant
	wire          sys_flash_tcm_chipselect_n_out_signal;                              // sys_flash:tcm_chipselect_n_out -> sys_flash_bridge:tcs_tcm_chipselect_n_out
	wire   [23:0] sys_flash_tcm_address_out_signal;                                   // sys_flash:tcm_address_out -> sys_flash_bridge:tcs_tcm_address_out
	wire   [31:0] sys_flash_tcm_data_out_signal;                                      // sys_flash:tcm_data_out -> sys_flash_bridge:tcs_tcm_data_out
	wire   [31:0] sys_flash_tcm_data_in;                                              // sys_flash_bridge:tcs_tcm_data_in -> sys_flash:tcm_data_in
	wire   [31:0] sys_cpu_data_master_readdata;                                       // mm_interconnect_0:sys_cpu_data_master_readdata -> sys_cpu:d_readdata
	wire          sys_cpu_data_master_waitrequest;                                    // mm_interconnect_0:sys_cpu_data_master_waitrequest -> sys_cpu:d_waitrequest
	wire          sys_cpu_data_master_debugaccess;                                    // sys_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:sys_cpu_data_master_debugaccess
	wire   [28:0] sys_cpu_data_master_address;                                        // sys_cpu:d_address -> mm_interconnect_0:sys_cpu_data_master_address
	wire    [3:0] sys_cpu_data_master_byteenable;                                     // sys_cpu:d_byteenable -> mm_interconnect_0:sys_cpu_data_master_byteenable
	wire          sys_cpu_data_master_read;                                           // sys_cpu:d_read -> mm_interconnect_0:sys_cpu_data_master_read
	wire          sys_cpu_data_master_readdatavalid;                                  // mm_interconnect_0:sys_cpu_data_master_readdatavalid -> sys_cpu:d_readdatavalid
	wire          sys_cpu_data_master_write;                                          // sys_cpu:d_write -> mm_interconnect_0:sys_cpu_data_master_write
	wire   [31:0] sys_cpu_data_master_writedata;                                      // sys_cpu:d_writedata -> mm_interconnect_0:sys_cpu_data_master_writedata
	wire   [31:0] sys_cpu_instruction_master_readdata;                                // mm_interconnect_0:sys_cpu_instruction_master_readdata -> sys_cpu:i_readdata
	wire          sys_cpu_instruction_master_waitrequest;                             // mm_interconnect_0:sys_cpu_instruction_master_waitrequest -> sys_cpu:i_waitrequest
	wire   [28:0] sys_cpu_instruction_master_address;                                 // sys_cpu:i_address -> mm_interconnect_0:sys_cpu_instruction_master_address
	wire          sys_cpu_instruction_master_read;                                    // sys_cpu:i_read -> mm_interconnect_0:sys_cpu_instruction_master_read
	wire          sys_cpu_instruction_master_readdatavalid;                           // mm_interconnect_0:sys_cpu_instruction_master_readdatavalid -> sys_cpu:i_readdatavalid
	wire    [1:0] axi_ad9680_dma_m_dest_axi_awburst;                                  // axi_ad9680_dma:m_dest_axi_awburst -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_awburst
	wire    [3:0] axi_ad9680_dma_m_dest_axi_arlen;                                    // axi_ad9680_dma:m_dest_axi_arlen -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_arlen
	wire   [15:0] axi_ad9680_dma_m_dest_axi_wstrb;                                    // axi_ad9680_dma:m_dest_axi_wstrb -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_wstrb
	wire          axi_ad9680_dma_m_dest_axi_wready;                                   // mm_interconnect_0:axi_ad9680_dma_m_dest_axi_wready -> axi_ad9680_dma:m_dest_axi_wready
	wire          axi_ad9680_dma_m_dest_axi_rid;                                      // mm_interconnect_0:axi_ad9680_dma_m_dest_axi_rid -> axi_ad9680_dma:m_dest_axi_rid
	wire          axi_ad9680_dma_m_dest_axi_rready;                                   // axi_ad9680_dma:m_dest_axi_rready -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_rready
	wire    [3:0] axi_ad9680_dma_m_dest_axi_awlen;                                    // axi_ad9680_dma:m_dest_axi_awlen -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_awlen
	wire          axi_ad9680_dma_m_dest_axi_wid;                                      // axi_ad9680_dma:m_dest_axi_wid -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_wid
	wire    [3:0] axi_ad9680_dma_m_dest_axi_arcache;                                  // axi_ad9680_dma:m_dest_axi_arcache -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_arcache
	wire          axi_ad9680_dma_m_dest_axi_wvalid;                                   // axi_ad9680_dma:m_dest_axi_wvalid -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_wvalid
	wire   [31:0] axi_ad9680_dma_m_dest_axi_araddr;                                   // axi_ad9680_dma:m_dest_axi_araddr -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_araddr
	wire    [2:0] axi_ad9680_dma_m_dest_axi_arprot;                                   // axi_ad9680_dma:m_dest_axi_arprot -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_arprot
	wire  [127:0] axi_ad9680_dma_m_dest_axi_wdata;                                    // axi_ad9680_dma:m_dest_axi_wdata -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_wdata
	wire          axi_ad9680_dma_m_dest_axi_arvalid;                                  // axi_ad9680_dma:m_dest_axi_arvalid -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_arvalid
	wire    [2:0] axi_ad9680_dma_m_dest_axi_awprot;                                   // axi_ad9680_dma:m_dest_axi_awprot -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_awprot
	wire    [3:0] axi_ad9680_dma_m_dest_axi_awcache;                                  // axi_ad9680_dma:m_dest_axi_awcache -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_awcache
	wire          axi_ad9680_dma_m_dest_axi_arid;                                     // axi_ad9680_dma:m_dest_axi_arid -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_arid
	wire    [1:0] axi_ad9680_dma_m_dest_axi_arlock;                                   // axi_ad9680_dma:m_dest_axi_arlock -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_arlock
	wire    [1:0] axi_ad9680_dma_m_dest_axi_awlock;                                   // axi_ad9680_dma:m_dest_axi_awlock -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_awlock
	wire   [31:0] axi_ad9680_dma_m_dest_axi_awaddr;                                   // axi_ad9680_dma:m_dest_axi_awaddr -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_awaddr
	wire    [1:0] axi_ad9680_dma_m_dest_axi_bresp;                                    // mm_interconnect_0:axi_ad9680_dma_m_dest_axi_bresp -> axi_ad9680_dma:m_dest_axi_bresp
	wire          axi_ad9680_dma_m_dest_axi_arready;                                  // mm_interconnect_0:axi_ad9680_dma_m_dest_axi_arready -> axi_ad9680_dma:m_dest_axi_arready
	wire  [127:0] axi_ad9680_dma_m_dest_axi_rdata;                                    // mm_interconnect_0:axi_ad9680_dma_m_dest_axi_rdata -> axi_ad9680_dma:m_dest_axi_rdata
	wire          axi_ad9680_dma_m_dest_axi_awready;                                  // mm_interconnect_0:axi_ad9680_dma_m_dest_axi_awready -> axi_ad9680_dma:m_dest_axi_awready
	wire    [1:0] axi_ad9680_dma_m_dest_axi_arburst;                                  // axi_ad9680_dma:m_dest_axi_arburst -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_arburst
	wire    [2:0] axi_ad9680_dma_m_dest_axi_arsize;                                   // axi_ad9680_dma:m_dest_axi_arsize -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_arsize
	wire          axi_ad9680_dma_m_dest_axi_bready;                                   // axi_ad9680_dma:m_dest_axi_bready -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_bready
	wire          axi_ad9680_dma_m_dest_axi_rlast;                                    // mm_interconnect_0:axi_ad9680_dma_m_dest_axi_rlast -> axi_ad9680_dma:m_dest_axi_rlast
	wire          axi_ad9680_dma_m_dest_axi_wlast;                                    // axi_ad9680_dma:m_dest_axi_wlast -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_wlast
	wire    [1:0] axi_ad9680_dma_m_dest_axi_rresp;                                    // mm_interconnect_0:axi_ad9680_dma_m_dest_axi_rresp -> axi_ad9680_dma:m_dest_axi_rresp
	wire          axi_ad9680_dma_m_dest_axi_awid;                                     // axi_ad9680_dma:m_dest_axi_awid -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_awid
	wire          axi_ad9680_dma_m_dest_axi_bid;                                      // mm_interconnect_0:axi_ad9680_dma_m_dest_axi_bid -> axi_ad9680_dma:m_dest_axi_bid
	wire          axi_ad9680_dma_m_dest_axi_bvalid;                                   // mm_interconnect_0:axi_ad9680_dma_m_dest_axi_bvalid -> axi_ad9680_dma:m_dest_axi_bvalid
	wire          axi_ad9680_dma_m_dest_axi_awvalid;                                  // axi_ad9680_dma:m_dest_axi_awvalid -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_awvalid
	wire          axi_ad9680_dma_m_dest_axi_rvalid;                                   // mm_interconnect_0:axi_ad9680_dma_m_dest_axi_rvalid -> axi_ad9680_dma:m_dest_axi_rvalid
	wire    [2:0] axi_ad9680_dma_m_dest_axi_awsize;                                   // axi_ad9680_dma:m_dest_axi_awsize -> mm_interconnect_0:axi_ad9680_dma_m_dest_axi_awsize
	wire    [1:0] axi_ad9144_dma_m_src_axi_awburst;                                   // axi_ad9144_dma:m_src_axi_awburst -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_awburst
	wire    [3:0] axi_ad9144_dma_m_src_axi_arlen;                                     // axi_ad9144_dma:m_src_axi_arlen -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_arlen
	wire   [15:0] axi_ad9144_dma_m_src_axi_wstrb;                                     // axi_ad9144_dma:m_src_axi_wstrb -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_wstrb
	wire          axi_ad9144_dma_m_src_axi_wready;                                    // mm_interconnect_0:axi_ad9144_dma_m_src_axi_wready -> axi_ad9144_dma:m_src_axi_wready
	wire          axi_ad9144_dma_m_src_axi_rid;                                       // mm_interconnect_0:axi_ad9144_dma_m_src_axi_rid -> axi_ad9144_dma:m_src_axi_rid
	wire          axi_ad9144_dma_m_src_axi_rready;                                    // axi_ad9144_dma:m_src_axi_rready -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_rready
	wire    [3:0] axi_ad9144_dma_m_src_axi_awlen;                                     // axi_ad9144_dma:m_src_axi_awlen -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_awlen
	wire          axi_ad9144_dma_m_src_axi_wid;                                       // axi_ad9144_dma:m_src_axi_wid -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_wid
	wire    [3:0] axi_ad9144_dma_m_src_axi_arcache;                                   // axi_ad9144_dma:m_src_axi_arcache -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_arcache
	wire          axi_ad9144_dma_m_src_axi_wvalid;                                    // axi_ad9144_dma:m_src_axi_wvalid -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_wvalid
	wire   [31:0] axi_ad9144_dma_m_src_axi_araddr;                                    // axi_ad9144_dma:m_src_axi_araddr -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_araddr
	wire    [2:0] axi_ad9144_dma_m_src_axi_arprot;                                    // axi_ad9144_dma:m_src_axi_arprot -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_arprot
	wire  [127:0] axi_ad9144_dma_m_src_axi_wdata;                                     // axi_ad9144_dma:m_src_axi_wdata -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_wdata
	wire          axi_ad9144_dma_m_src_axi_arvalid;                                   // axi_ad9144_dma:m_src_axi_arvalid -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_arvalid
	wire    [2:0] axi_ad9144_dma_m_src_axi_awprot;                                    // axi_ad9144_dma:m_src_axi_awprot -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_awprot
	wire    [3:0] axi_ad9144_dma_m_src_axi_awcache;                                   // axi_ad9144_dma:m_src_axi_awcache -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_awcache
	wire          axi_ad9144_dma_m_src_axi_arid;                                      // axi_ad9144_dma:m_src_axi_arid -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_arid
	wire    [1:0] axi_ad9144_dma_m_src_axi_arlock;                                    // axi_ad9144_dma:m_src_axi_arlock -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_arlock
	wire    [1:0] axi_ad9144_dma_m_src_axi_awlock;                                    // axi_ad9144_dma:m_src_axi_awlock -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_awlock
	wire   [31:0] axi_ad9144_dma_m_src_axi_awaddr;                                    // axi_ad9144_dma:m_src_axi_awaddr -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_awaddr
	wire    [1:0] axi_ad9144_dma_m_src_axi_bresp;                                     // mm_interconnect_0:axi_ad9144_dma_m_src_axi_bresp -> axi_ad9144_dma:m_src_axi_bresp
	wire          axi_ad9144_dma_m_src_axi_arready;                                   // mm_interconnect_0:axi_ad9144_dma_m_src_axi_arready -> axi_ad9144_dma:m_src_axi_arready
	wire  [127:0] axi_ad9144_dma_m_src_axi_rdata;                                     // mm_interconnect_0:axi_ad9144_dma_m_src_axi_rdata -> axi_ad9144_dma:m_src_axi_rdata
	wire          axi_ad9144_dma_m_src_axi_awready;                                   // mm_interconnect_0:axi_ad9144_dma_m_src_axi_awready -> axi_ad9144_dma:m_src_axi_awready
	wire    [1:0] axi_ad9144_dma_m_src_axi_arburst;                                   // axi_ad9144_dma:m_src_axi_arburst -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_arburst
	wire    [2:0] axi_ad9144_dma_m_src_axi_arsize;                                    // axi_ad9144_dma:m_src_axi_arsize -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_arsize
	wire          axi_ad9144_dma_m_src_axi_bready;                                    // axi_ad9144_dma:m_src_axi_bready -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_bready
	wire          axi_ad9144_dma_m_src_axi_rlast;                                     // mm_interconnect_0:axi_ad9144_dma_m_src_axi_rlast -> axi_ad9144_dma:m_src_axi_rlast
	wire          axi_ad9144_dma_m_src_axi_wlast;                                     // axi_ad9144_dma:m_src_axi_wlast -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_wlast
	wire    [1:0] axi_ad9144_dma_m_src_axi_rresp;                                     // mm_interconnect_0:axi_ad9144_dma_m_src_axi_rresp -> axi_ad9144_dma:m_src_axi_rresp
	wire          axi_ad9144_dma_m_src_axi_awid;                                      // axi_ad9144_dma:m_src_axi_awid -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_awid
	wire          axi_ad9144_dma_m_src_axi_bid;                                       // mm_interconnect_0:axi_ad9144_dma_m_src_axi_bid -> axi_ad9144_dma:m_src_axi_bid
	wire          axi_ad9144_dma_m_src_axi_bvalid;                                    // mm_interconnect_0:axi_ad9144_dma_m_src_axi_bvalid -> axi_ad9144_dma:m_src_axi_bvalid
	wire          axi_ad9144_dma_m_src_axi_awvalid;                                   // axi_ad9144_dma:m_src_axi_awvalid -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_awvalid
	wire          axi_ad9144_dma_m_src_axi_rvalid;                                    // mm_interconnect_0:axi_ad9144_dma_m_src_axi_rvalid -> axi_ad9144_dma:m_src_axi_rvalid
	wire    [2:0] axi_ad9144_dma_m_src_axi_awsize;                                    // axi_ad9144_dma:m_src_axi_awsize -> mm_interconnect_0:axi_ad9144_dma_m_src_axi_awsize
	wire   [63:0] sys_ethernet_dma_tx_mm_read_readdata;                               // mm_interconnect_0:sys_ethernet_dma_tx_mm_read_readdata -> sys_ethernet_dma_tx:mm_read_readdata
	wire          sys_ethernet_dma_tx_mm_read_waitrequest;                            // mm_interconnect_0:sys_ethernet_dma_tx_mm_read_waitrequest -> sys_ethernet_dma_tx:mm_read_waitrequest
	wire   [31:0] sys_ethernet_dma_tx_mm_read_address;                                // sys_ethernet_dma_tx:mm_read_address -> mm_interconnect_0:sys_ethernet_dma_tx_mm_read_address
	wire          sys_ethernet_dma_tx_mm_read_read;                                   // sys_ethernet_dma_tx:mm_read_read -> mm_interconnect_0:sys_ethernet_dma_tx_mm_read_read
	wire    [7:0] sys_ethernet_dma_tx_mm_read_byteenable;                             // sys_ethernet_dma_tx:mm_read_byteenable -> mm_interconnect_0:sys_ethernet_dma_tx_mm_read_byteenable
	wire          sys_ethernet_dma_tx_mm_read_readdatavalid;                          // mm_interconnect_0:sys_ethernet_dma_tx_mm_read_readdatavalid -> sys_ethernet_dma_tx:mm_read_readdatavalid
	wire    [6:0] sys_ethernet_dma_tx_mm_read_burstcount;                             // sys_ethernet_dma_tx:mm_read_burstcount -> mm_interconnect_0:sys_ethernet_dma_tx_mm_read_burstcount
	wire          sys_ethernet_dma_rx_mm_write_waitrequest;                           // mm_interconnect_0:sys_ethernet_dma_rx_mm_write_waitrequest -> sys_ethernet_dma_rx:mm_write_waitrequest
	wire   [31:0] sys_ethernet_dma_rx_mm_write_address;                               // sys_ethernet_dma_rx:mm_write_address -> mm_interconnect_0:sys_ethernet_dma_rx_mm_write_address
	wire    [7:0] sys_ethernet_dma_rx_mm_write_byteenable;                            // sys_ethernet_dma_rx:mm_write_byteenable -> mm_interconnect_0:sys_ethernet_dma_rx_mm_write_byteenable
	wire          sys_ethernet_dma_rx_mm_write_write;                                 // sys_ethernet_dma_rx:mm_write_write -> mm_interconnect_0:sys_ethernet_dma_rx_mm_write_write
	wire   [63:0] sys_ethernet_dma_rx_mm_write_writedata;                             // sys_ethernet_dma_rx:mm_write_writedata -> mm_interconnect_0:sys_ethernet_dma_rx_mm_write_writedata
	wire    [6:0] sys_ethernet_dma_rx_mm_write_burstcount;                            // sys_ethernet_dma_rx:mm_write_burstcount -> mm_interconnect_0:sys_ethernet_dma_rx_mm_write_burstcount
	wire          mm_interconnect_0_sys_uart_avalon_jtag_slave_chipselect;            // mm_interconnect_0:sys_uart_avalon_jtag_slave_chipselect -> sys_uart:av_chipselect
	wire   [31:0] mm_interconnect_0_sys_uart_avalon_jtag_slave_readdata;              // sys_uart:av_readdata -> mm_interconnect_0:sys_uart_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_sys_uart_avalon_jtag_slave_waitrequest;           // sys_uart:av_waitrequest -> mm_interconnect_0:sys_uart_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_sys_uart_avalon_jtag_slave_address;               // mm_interconnect_0:sys_uart_avalon_jtag_slave_address -> sys_uart:av_address
	wire          mm_interconnect_0_sys_uart_avalon_jtag_slave_read;                  // mm_interconnect_0:sys_uart_avalon_jtag_slave_read -> sys_uart:av_read_n
	wire          mm_interconnect_0_sys_uart_avalon_jtag_slave_write;                 // mm_interconnect_0:sys_uart_avalon_jtag_slave_write -> sys_uart:av_write_n
	wire   [31:0] mm_interconnect_0_sys_uart_avalon_jtag_slave_writedata;             // mm_interconnect_0:sys_uart_avalon_jtag_slave_writedata -> sys_uart:av_writedata
	wire   [31:0] mm_interconnect_0_sys_ethernet_control_port_readdata;               // sys_ethernet:reg_data_out -> mm_interconnect_0:sys_ethernet_control_port_readdata
	wire          mm_interconnect_0_sys_ethernet_control_port_waitrequest;            // sys_ethernet:reg_busy -> mm_interconnect_0:sys_ethernet_control_port_waitrequest
	wire    [7:0] mm_interconnect_0_sys_ethernet_control_port_address;                // mm_interconnect_0:sys_ethernet_control_port_address -> sys_ethernet:reg_addr
	wire          mm_interconnect_0_sys_ethernet_control_port_read;                   // mm_interconnect_0:sys_ethernet_control_port_read -> sys_ethernet:reg_rd
	wire          mm_interconnect_0_sys_ethernet_control_port_write;                  // mm_interconnect_0:sys_ethernet_control_port_write -> sys_ethernet:reg_wr
	wire   [31:0] mm_interconnect_0_sys_ethernet_control_port_writedata;              // mm_interconnect_0:sys_ethernet_control_port_writedata -> sys_ethernet:reg_data_in
	wire   [31:0] mm_interconnect_0_sys_id_control_slave_readdata;                    // sys_id:readdata -> mm_interconnect_0:sys_id_control_slave_readdata
	wire    [0:0] mm_interconnect_0_sys_id_control_slave_address;                     // mm_interconnect_0:sys_id_control_slave_address -> sys_id:address
	wire   [31:0] mm_interconnect_0_sys_ethernet_dma_rx_csr_readdata;                 // sys_ethernet_dma_rx:csr_readdata -> mm_interconnect_0:sys_ethernet_dma_rx_csr_readdata
	wire    [2:0] mm_interconnect_0_sys_ethernet_dma_rx_csr_address;                  // mm_interconnect_0:sys_ethernet_dma_rx_csr_address -> sys_ethernet_dma_rx:csr_address
	wire          mm_interconnect_0_sys_ethernet_dma_rx_csr_read;                     // mm_interconnect_0:sys_ethernet_dma_rx_csr_read -> sys_ethernet_dma_rx:csr_read
	wire    [3:0] mm_interconnect_0_sys_ethernet_dma_rx_csr_byteenable;               // mm_interconnect_0:sys_ethernet_dma_rx_csr_byteenable -> sys_ethernet_dma_rx:csr_byteenable
	wire          mm_interconnect_0_sys_ethernet_dma_rx_csr_write;                    // mm_interconnect_0:sys_ethernet_dma_rx_csr_write -> sys_ethernet_dma_rx:csr_write
	wire   [31:0] mm_interconnect_0_sys_ethernet_dma_rx_csr_writedata;                // mm_interconnect_0:sys_ethernet_dma_rx_csr_writedata -> sys_ethernet_dma_rx:csr_writedata
	wire   [31:0] mm_interconnect_0_sys_ethernet_dma_tx_csr_readdata;                 // sys_ethernet_dma_tx:csr_readdata -> mm_interconnect_0:sys_ethernet_dma_tx_csr_readdata
	wire    [2:0] mm_interconnect_0_sys_ethernet_dma_tx_csr_address;                  // mm_interconnect_0:sys_ethernet_dma_tx_csr_address -> sys_ethernet_dma_tx:csr_address
	wire          mm_interconnect_0_sys_ethernet_dma_tx_csr_read;                     // mm_interconnect_0:sys_ethernet_dma_tx_csr_read -> sys_ethernet_dma_tx:csr_read
	wire    [3:0] mm_interconnect_0_sys_ethernet_dma_tx_csr_byteenable;               // mm_interconnect_0:sys_ethernet_dma_tx_csr_byteenable -> sys_ethernet_dma_tx:csr_byteenable
	wire          mm_interconnect_0_sys_ethernet_dma_tx_csr_write;                    // mm_interconnect_0:sys_ethernet_dma_tx_csr_write -> sys_ethernet_dma_tx:csr_write
	wire   [31:0] mm_interconnect_0_sys_ethernet_dma_tx_csr_writedata;                // mm_interconnect_0:sys_ethernet_dma_tx_csr_writedata -> sys_ethernet_dma_tx:csr_writedata
	wire  [511:0] mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_readdata;               // sys_ddr3_cntrl:amm_readdata_0 -> mm_interconnect_0:sys_ddr3_cntrl_ctrl_amm_0_readdata
	wire          mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_waitrequest;            // sys_ddr3_cntrl:amm_ready_0 -> mm_interconnect_0:sys_ddr3_cntrl_ctrl_amm_0_waitrequest
	wire   [21:0] mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_address;                // mm_interconnect_0:sys_ddr3_cntrl_ctrl_amm_0_address -> sys_ddr3_cntrl:amm_address_0
	wire          mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_read;                   // mm_interconnect_0:sys_ddr3_cntrl_ctrl_amm_0_read -> sys_ddr3_cntrl:amm_read_0
	wire   [63:0] mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_byteenable;             // mm_interconnect_0:sys_ddr3_cntrl_ctrl_amm_0_byteenable -> sys_ddr3_cntrl:amm_byteenable_0
	wire          mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_readdatavalid;          // sys_ddr3_cntrl:amm_readdatavalid_0 -> mm_interconnect_0:sys_ddr3_cntrl_ctrl_amm_0_readdatavalid
	wire          mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_write;                  // mm_interconnect_0:sys_ddr3_cntrl_ctrl_amm_0_write -> sys_ddr3_cntrl:amm_write_0
	wire  [511:0] mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_writedata;              // mm_interconnect_0:sys_ddr3_cntrl_ctrl_amm_0_writedata -> sys_ddr3_cntrl:amm_writedata_0
	wire    [6:0] mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_burstcount;             // mm_interconnect_0:sys_ddr3_cntrl_ctrl_amm_0_burstcount -> sys_ddr3_cntrl:amm_burstcount_0
	wire   [31:0] mm_interconnect_0_sys_cpu_debug_mem_slave_readdata;                 // sys_cpu:debug_mem_slave_readdata -> mm_interconnect_0:sys_cpu_debug_mem_slave_readdata
	wire          mm_interconnect_0_sys_cpu_debug_mem_slave_waitrequest;              // sys_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:sys_cpu_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_sys_cpu_debug_mem_slave_debugaccess;              // mm_interconnect_0:sys_cpu_debug_mem_slave_debugaccess -> sys_cpu:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_sys_cpu_debug_mem_slave_address;                  // mm_interconnect_0:sys_cpu_debug_mem_slave_address -> sys_cpu:debug_mem_slave_address
	wire          mm_interconnect_0_sys_cpu_debug_mem_slave_read;                     // mm_interconnect_0:sys_cpu_debug_mem_slave_read -> sys_cpu:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_sys_cpu_debug_mem_slave_byteenable;               // mm_interconnect_0:sys_cpu_debug_mem_slave_byteenable -> sys_cpu:debug_mem_slave_byteenable
	wire          mm_interconnect_0_sys_cpu_debug_mem_slave_write;                    // mm_interconnect_0:sys_cpu_debug_mem_slave_write -> sys_cpu:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_sys_cpu_debug_mem_slave_writedata;                // mm_interconnect_0:sys_cpu_debug_mem_slave_writedata -> sys_cpu:debug_mem_slave_writedata
	wire          mm_interconnect_0_sys_ethernet_dma_rx_descriptor_slave_waitrequest; // sys_ethernet_dma_rx:descriptor_slave_waitrequest -> mm_interconnect_0:sys_ethernet_dma_rx_descriptor_slave_waitrequest
	wire   [31:0] mm_interconnect_0_sys_ethernet_dma_rx_descriptor_slave_byteenable;  // mm_interconnect_0:sys_ethernet_dma_rx_descriptor_slave_byteenable -> sys_ethernet_dma_rx:descriptor_slave_byteenable
	wire          mm_interconnect_0_sys_ethernet_dma_rx_descriptor_slave_write;       // mm_interconnect_0:sys_ethernet_dma_rx_descriptor_slave_write -> sys_ethernet_dma_rx:descriptor_slave_write
	wire  [255:0] mm_interconnect_0_sys_ethernet_dma_rx_descriptor_slave_writedata;   // mm_interconnect_0:sys_ethernet_dma_rx_descriptor_slave_writedata -> sys_ethernet_dma_rx:descriptor_slave_writedata
	wire          mm_interconnect_0_sys_ethernet_dma_tx_descriptor_slave_waitrequest; // sys_ethernet_dma_tx:descriptor_slave_waitrequest -> mm_interconnect_0:sys_ethernet_dma_tx_descriptor_slave_waitrequest
	wire   [31:0] mm_interconnect_0_sys_ethernet_dma_tx_descriptor_slave_byteenable;  // mm_interconnect_0:sys_ethernet_dma_tx_descriptor_slave_byteenable -> sys_ethernet_dma_tx:descriptor_slave_byteenable
	wire          mm_interconnect_0_sys_ethernet_dma_tx_descriptor_slave_write;       // mm_interconnect_0:sys_ethernet_dma_tx_descriptor_slave_write -> sys_ethernet_dma_tx:descriptor_slave_write
	wire  [255:0] mm_interconnect_0_sys_ethernet_dma_tx_descriptor_slave_writedata;   // mm_interconnect_0:sys_ethernet_dma_tx_descriptor_slave_writedata -> sys_ethernet_dma_tx:descriptor_slave_writedata
	wire   [31:0] mm_interconnect_0_avl_adxcfg_0_rcfg_s0_readdata;                    // avl_adxcfg_0:rcfg_in_readdata_0 -> mm_interconnect_0:avl_adxcfg_0_rcfg_s0_readdata
	wire          mm_interconnect_0_avl_adxcfg_0_rcfg_s0_waitrequest;                 // avl_adxcfg_0:rcfg_in_waitrequest_0 -> mm_interconnect_0:avl_adxcfg_0_rcfg_s0_waitrequest
	wire    [9:0] mm_interconnect_0_avl_adxcfg_0_rcfg_s0_address;                     // mm_interconnect_0:avl_adxcfg_0_rcfg_s0_address -> avl_adxcfg_0:rcfg_in_address_0
	wire          mm_interconnect_0_avl_adxcfg_0_rcfg_s0_read;                        // mm_interconnect_0:avl_adxcfg_0_rcfg_s0_read -> avl_adxcfg_0:rcfg_in_read_0
	wire          mm_interconnect_0_avl_adxcfg_0_rcfg_s0_write;                       // mm_interconnect_0:avl_adxcfg_0_rcfg_s0_write -> avl_adxcfg_0:rcfg_in_write_0
	wire   [31:0] mm_interconnect_0_avl_adxcfg_0_rcfg_s0_writedata;                   // mm_interconnect_0:avl_adxcfg_0_rcfg_s0_writedata -> avl_adxcfg_0:rcfg_in_writedata_0
	wire   [31:0] mm_interconnect_0_avl_adxcfg_1_rcfg_s0_readdata;                    // avl_adxcfg_1:rcfg_in_readdata_0 -> mm_interconnect_0:avl_adxcfg_1_rcfg_s0_readdata
	wire          mm_interconnect_0_avl_adxcfg_1_rcfg_s0_waitrequest;                 // avl_adxcfg_1:rcfg_in_waitrequest_0 -> mm_interconnect_0:avl_adxcfg_1_rcfg_s0_waitrequest
	wire    [9:0] mm_interconnect_0_avl_adxcfg_1_rcfg_s0_address;                     // mm_interconnect_0:avl_adxcfg_1_rcfg_s0_address -> avl_adxcfg_1:rcfg_in_address_0
	wire          mm_interconnect_0_avl_adxcfg_1_rcfg_s0_read;                        // mm_interconnect_0:avl_adxcfg_1_rcfg_s0_read -> avl_adxcfg_1:rcfg_in_read_0
	wire          mm_interconnect_0_avl_adxcfg_1_rcfg_s0_write;                       // mm_interconnect_0:avl_adxcfg_1_rcfg_s0_write -> avl_adxcfg_1:rcfg_in_write_0
	wire   [31:0] mm_interconnect_0_avl_adxcfg_1_rcfg_s0_writedata;                   // mm_interconnect_0:avl_adxcfg_1_rcfg_s0_writedata -> avl_adxcfg_1:rcfg_in_writedata_0
	wire   [31:0] mm_interconnect_0_avl_adxcfg_2_rcfg_s0_readdata;                    // avl_adxcfg_2:rcfg_in_readdata_0 -> mm_interconnect_0:avl_adxcfg_2_rcfg_s0_readdata
	wire          mm_interconnect_0_avl_adxcfg_2_rcfg_s0_waitrequest;                 // avl_adxcfg_2:rcfg_in_waitrequest_0 -> mm_interconnect_0:avl_adxcfg_2_rcfg_s0_waitrequest
	wire    [9:0] mm_interconnect_0_avl_adxcfg_2_rcfg_s0_address;                     // mm_interconnect_0:avl_adxcfg_2_rcfg_s0_address -> avl_adxcfg_2:rcfg_in_address_0
	wire          mm_interconnect_0_avl_adxcfg_2_rcfg_s0_read;                        // mm_interconnect_0:avl_adxcfg_2_rcfg_s0_read -> avl_adxcfg_2:rcfg_in_read_0
	wire          mm_interconnect_0_avl_adxcfg_2_rcfg_s0_write;                       // mm_interconnect_0:avl_adxcfg_2_rcfg_s0_write -> avl_adxcfg_2:rcfg_in_write_0
	wire   [31:0] mm_interconnect_0_avl_adxcfg_2_rcfg_s0_writedata;                   // mm_interconnect_0:avl_adxcfg_2_rcfg_s0_writedata -> avl_adxcfg_2:rcfg_in_writedata_0
	wire   [31:0] mm_interconnect_0_avl_adxcfg_3_rcfg_s0_readdata;                    // avl_adxcfg_3:rcfg_in_readdata_0 -> mm_interconnect_0:avl_adxcfg_3_rcfg_s0_readdata
	wire          mm_interconnect_0_avl_adxcfg_3_rcfg_s0_waitrequest;                 // avl_adxcfg_3:rcfg_in_waitrequest_0 -> mm_interconnect_0:avl_adxcfg_3_rcfg_s0_waitrequest
	wire    [9:0] mm_interconnect_0_avl_adxcfg_3_rcfg_s0_address;                     // mm_interconnect_0:avl_adxcfg_3_rcfg_s0_address -> avl_adxcfg_3:rcfg_in_address_0
	wire          mm_interconnect_0_avl_adxcfg_3_rcfg_s0_read;                        // mm_interconnect_0:avl_adxcfg_3_rcfg_s0_read -> avl_adxcfg_3:rcfg_in_read_0
	wire          mm_interconnect_0_avl_adxcfg_3_rcfg_s0_write;                       // mm_interconnect_0:avl_adxcfg_3_rcfg_s0_write -> avl_adxcfg_3:rcfg_in_write_0
	wire   [31:0] mm_interconnect_0_avl_adxcfg_3_rcfg_s0_writedata;                   // mm_interconnect_0:avl_adxcfg_3_rcfg_s0_writedata -> avl_adxcfg_3:rcfg_in_writedata_0
	wire   [31:0] mm_interconnect_0_avl_adxcfg_0_rcfg_s1_readdata;                    // avl_adxcfg_0:rcfg_in_readdata_1 -> mm_interconnect_0:avl_adxcfg_0_rcfg_s1_readdata
	wire          mm_interconnect_0_avl_adxcfg_0_rcfg_s1_waitrequest;                 // avl_adxcfg_0:rcfg_in_waitrequest_1 -> mm_interconnect_0:avl_adxcfg_0_rcfg_s1_waitrequest
	wire    [9:0] mm_interconnect_0_avl_adxcfg_0_rcfg_s1_address;                     // mm_interconnect_0:avl_adxcfg_0_rcfg_s1_address -> avl_adxcfg_0:rcfg_in_address_1
	wire          mm_interconnect_0_avl_adxcfg_0_rcfg_s1_read;                        // mm_interconnect_0:avl_adxcfg_0_rcfg_s1_read -> avl_adxcfg_0:rcfg_in_read_1
	wire          mm_interconnect_0_avl_adxcfg_0_rcfg_s1_write;                       // mm_interconnect_0:avl_adxcfg_0_rcfg_s1_write -> avl_adxcfg_0:rcfg_in_write_1
	wire   [31:0] mm_interconnect_0_avl_adxcfg_0_rcfg_s1_writedata;                   // mm_interconnect_0:avl_adxcfg_0_rcfg_s1_writedata -> avl_adxcfg_0:rcfg_in_writedata_1
	wire   [31:0] mm_interconnect_0_avl_adxcfg_1_rcfg_s1_readdata;                    // avl_adxcfg_1:rcfg_in_readdata_1 -> mm_interconnect_0:avl_adxcfg_1_rcfg_s1_readdata
	wire          mm_interconnect_0_avl_adxcfg_1_rcfg_s1_waitrequest;                 // avl_adxcfg_1:rcfg_in_waitrequest_1 -> mm_interconnect_0:avl_adxcfg_1_rcfg_s1_waitrequest
	wire    [9:0] mm_interconnect_0_avl_adxcfg_1_rcfg_s1_address;                     // mm_interconnect_0:avl_adxcfg_1_rcfg_s1_address -> avl_adxcfg_1:rcfg_in_address_1
	wire          mm_interconnect_0_avl_adxcfg_1_rcfg_s1_read;                        // mm_interconnect_0:avl_adxcfg_1_rcfg_s1_read -> avl_adxcfg_1:rcfg_in_read_1
	wire          mm_interconnect_0_avl_adxcfg_1_rcfg_s1_write;                       // mm_interconnect_0:avl_adxcfg_1_rcfg_s1_write -> avl_adxcfg_1:rcfg_in_write_1
	wire   [31:0] mm_interconnect_0_avl_adxcfg_1_rcfg_s1_writedata;                   // mm_interconnect_0:avl_adxcfg_1_rcfg_s1_writedata -> avl_adxcfg_1:rcfg_in_writedata_1
	wire   [31:0] mm_interconnect_0_avl_adxcfg_2_rcfg_s1_readdata;                    // avl_adxcfg_2:rcfg_in_readdata_1 -> mm_interconnect_0:avl_adxcfg_2_rcfg_s1_readdata
	wire          mm_interconnect_0_avl_adxcfg_2_rcfg_s1_waitrequest;                 // avl_adxcfg_2:rcfg_in_waitrequest_1 -> mm_interconnect_0:avl_adxcfg_2_rcfg_s1_waitrequest
	wire    [9:0] mm_interconnect_0_avl_adxcfg_2_rcfg_s1_address;                     // mm_interconnect_0:avl_adxcfg_2_rcfg_s1_address -> avl_adxcfg_2:rcfg_in_address_1
	wire          mm_interconnect_0_avl_adxcfg_2_rcfg_s1_read;                        // mm_interconnect_0:avl_adxcfg_2_rcfg_s1_read -> avl_adxcfg_2:rcfg_in_read_1
	wire          mm_interconnect_0_avl_adxcfg_2_rcfg_s1_write;                       // mm_interconnect_0:avl_adxcfg_2_rcfg_s1_write -> avl_adxcfg_2:rcfg_in_write_1
	wire   [31:0] mm_interconnect_0_avl_adxcfg_2_rcfg_s1_writedata;                   // mm_interconnect_0:avl_adxcfg_2_rcfg_s1_writedata -> avl_adxcfg_2:rcfg_in_writedata_1
	wire   [31:0] mm_interconnect_0_avl_adxcfg_3_rcfg_s1_readdata;                    // avl_adxcfg_3:rcfg_in_readdata_1 -> mm_interconnect_0:avl_adxcfg_3_rcfg_s1_readdata
	wire          mm_interconnect_0_avl_adxcfg_3_rcfg_s1_waitrequest;                 // avl_adxcfg_3:rcfg_in_waitrequest_1 -> mm_interconnect_0:avl_adxcfg_3_rcfg_s1_waitrequest
	wire    [9:0] mm_interconnect_0_avl_adxcfg_3_rcfg_s1_address;                     // mm_interconnect_0:avl_adxcfg_3_rcfg_s1_address -> avl_adxcfg_3:rcfg_in_address_1
	wire          mm_interconnect_0_avl_adxcfg_3_rcfg_s1_read;                        // mm_interconnect_0:avl_adxcfg_3_rcfg_s1_read -> avl_adxcfg_3:rcfg_in_read_1
	wire          mm_interconnect_0_avl_adxcfg_3_rcfg_s1_write;                       // mm_interconnect_0:avl_adxcfg_3_rcfg_s1_write -> avl_adxcfg_3:rcfg_in_write_1
	wire   [31:0] mm_interconnect_0_avl_adxcfg_3_rcfg_s1_writedata;                   // mm_interconnect_0:avl_adxcfg_3_rcfg_s1_writedata -> avl_adxcfg_3:rcfg_in_writedata_1
	wire   [31:0] mm_interconnect_0_sys_ethernet_dma_rx_response_readdata;            // sys_ethernet_dma_rx:response_readdata -> mm_interconnect_0:sys_ethernet_dma_rx_response_readdata
	wire          mm_interconnect_0_sys_ethernet_dma_rx_response_waitrequest;         // sys_ethernet_dma_rx:response_waitrequest -> mm_interconnect_0:sys_ethernet_dma_rx_response_waitrequest
	wire    [0:0] mm_interconnect_0_sys_ethernet_dma_rx_response_address;             // mm_interconnect_0:sys_ethernet_dma_rx_response_address -> sys_ethernet_dma_rx:response_address
	wire          mm_interconnect_0_sys_ethernet_dma_rx_response_read;                // mm_interconnect_0:sys_ethernet_dma_rx_response_read -> sys_ethernet_dma_rx:response_read
	wire    [3:0] mm_interconnect_0_sys_ethernet_dma_rx_response_byteenable;          // mm_interconnect_0:sys_ethernet_dma_rx_response_byteenable -> sys_ethernet_dma_rx:response_byteenable
	wire          mm_interconnect_0_sys_int_mem_s1_chipselect;                        // mm_interconnect_0:sys_int_mem_s1_chipselect -> sys_int_mem:chipselect
	wire   [31:0] mm_interconnect_0_sys_int_mem_s1_readdata;                          // sys_int_mem:readdata -> mm_interconnect_0:sys_int_mem_s1_readdata
	wire   [15:0] mm_interconnect_0_sys_int_mem_s1_address;                           // mm_interconnect_0:sys_int_mem_s1_address -> sys_int_mem:address
	wire    [3:0] mm_interconnect_0_sys_int_mem_s1_byteenable;                        // mm_interconnect_0:sys_int_mem_s1_byteenable -> sys_int_mem:byteenable
	wire          mm_interconnect_0_sys_int_mem_s1_write;                             // mm_interconnect_0:sys_int_mem_s1_write -> sys_int_mem:write
	wire   [31:0] mm_interconnect_0_sys_int_mem_s1_writedata;                         // mm_interconnect_0:sys_int_mem_s1_writedata -> sys_int_mem:writedata
	wire          mm_interconnect_0_sys_int_mem_s1_clken;                             // mm_interconnect_0:sys_int_mem_s1_clken -> sys_int_mem:clken
	wire          mm_interconnect_0_sys_timer_1_s1_chipselect;                        // mm_interconnect_0:sys_timer_1_s1_chipselect -> sys_timer_1:chipselect
	wire   [15:0] mm_interconnect_0_sys_timer_1_s1_readdata;                          // sys_timer_1:readdata -> mm_interconnect_0:sys_timer_1_s1_readdata
	wire    [2:0] mm_interconnect_0_sys_timer_1_s1_address;                           // mm_interconnect_0:sys_timer_1_s1_address -> sys_timer_1:address
	wire          mm_interconnect_0_sys_timer_1_s1_write;                             // mm_interconnect_0:sys_timer_1_s1_write -> sys_timer_1:write_n
	wire   [15:0] mm_interconnect_0_sys_timer_1_s1_writedata;                         // mm_interconnect_0:sys_timer_1_s1_writedata -> sys_timer_1:writedata
	wire          mm_interconnect_0_sys_timer_2_s1_chipselect;                        // mm_interconnect_0:sys_timer_2_s1_chipselect -> sys_timer_2:chipselect
	wire   [15:0] mm_interconnect_0_sys_timer_2_s1_readdata;                          // sys_timer_2:readdata -> mm_interconnect_0:sys_timer_2_s1_readdata
	wire    [2:0] mm_interconnect_0_sys_timer_2_s1_address;                           // mm_interconnect_0:sys_timer_2_s1_address -> sys_timer_2:address
	wire          mm_interconnect_0_sys_timer_2_s1_write;                             // mm_interconnect_0:sys_timer_2_s1_write -> sys_timer_2:write_n
	wire   [15:0] mm_interconnect_0_sys_timer_2_s1_writedata;                         // mm_interconnect_0:sys_timer_2_s1_writedata -> sys_timer_2:writedata
	wire          mm_interconnect_0_sys_gpio_bd_s1_chipselect;                        // mm_interconnect_0:sys_gpio_bd_s1_chipselect -> sys_gpio_bd:chipselect
	wire   [31:0] mm_interconnect_0_sys_gpio_bd_s1_readdata;                          // sys_gpio_bd:readdata -> mm_interconnect_0:sys_gpio_bd_s1_readdata
	wire    [1:0] mm_interconnect_0_sys_gpio_bd_s1_address;                           // mm_interconnect_0:sys_gpio_bd_s1_address -> sys_gpio_bd:address
	wire          mm_interconnect_0_sys_gpio_bd_s1_write;                             // mm_interconnect_0:sys_gpio_bd_s1_write -> sys_gpio_bd:write_n
	wire   [31:0] mm_interconnect_0_sys_gpio_bd_s1_writedata;                         // mm_interconnect_0:sys_gpio_bd_s1_writedata -> sys_gpio_bd:writedata
	wire          mm_interconnect_0_sys_gpio_in_s1_chipselect;                        // mm_interconnect_0:sys_gpio_in_s1_chipselect -> sys_gpio_in:chipselect
	wire   [31:0] mm_interconnect_0_sys_gpio_in_s1_readdata;                          // sys_gpio_in:readdata -> mm_interconnect_0:sys_gpio_in_s1_readdata
	wire    [1:0] mm_interconnect_0_sys_gpio_in_s1_address;                           // mm_interconnect_0:sys_gpio_in_s1_address -> sys_gpio_in:address
	wire          mm_interconnect_0_sys_gpio_in_s1_write;                             // mm_interconnect_0:sys_gpio_in_s1_write -> sys_gpio_in:write_n
	wire   [31:0] mm_interconnect_0_sys_gpio_in_s1_writedata;                         // mm_interconnect_0:sys_gpio_in_s1_writedata -> sys_gpio_in:writedata
	wire          mm_interconnect_0_sys_gpio_out_s1_chipselect;                       // mm_interconnect_0:sys_gpio_out_s1_chipselect -> sys_gpio_out:chipselect
	wire   [31:0] mm_interconnect_0_sys_gpio_out_s1_readdata;                         // sys_gpio_out:readdata -> mm_interconnect_0:sys_gpio_out_s1_readdata
	wire    [1:0] mm_interconnect_0_sys_gpio_out_s1_address;                          // mm_interconnect_0:sys_gpio_out_s1_address -> sys_gpio_out:address
	wire          mm_interconnect_0_sys_gpio_out_s1_write;                            // mm_interconnect_0:sys_gpio_out_s1_write -> sys_gpio_out:write_n
	wire   [31:0] mm_interconnect_0_sys_gpio_out_s1_writedata;                        // mm_interconnect_0:sys_gpio_out_s1_writedata -> sys_gpio_out:writedata
	wire   [11:0] mm_interconnect_0_axi_ad9144_dma_s_axi_awaddr;                      // mm_interconnect_0:axi_ad9144_dma_s_axi_awaddr -> axi_ad9144_dma:s_axi_awaddr
	wire    [1:0] mm_interconnect_0_axi_ad9144_dma_s_axi_bresp;                       // axi_ad9144_dma:s_axi_bresp -> mm_interconnect_0:axi_ad9144_dma_s_axi_bresp
	wire          mm_interconnect_0_axi_ad9144_dma_s_axi_arready;                     // axi_ad9144_dma:s_axi_arready -> mm_interconnect_0:axi_ad9144_dma_s_axi_arready
	wire   [31:0] mm_interconnect_0_axi_ad9144_dma_s_axi_rdata;                       // axi_ad9144_dma:s_axi_rdata -> mm_interconnect_0:axi_ad9144_dma_s_axi_rdata
	wire    [3:0] mm_interconnect_0_axi_ad9144_dma_s_axi_wstrb;                       // mm_interconnect_0:axi_ad9144_dma_s_axi_wstrb -> axi_ad9144_dma:s_axi_wstrb
	wire          mm_interconnect_0_axi_ad9144_dma_s_axi_wready;                      // axi_ad9144_dma:s_axi_wready -> mm_interconnect_0:axi_ad9144_dma_s_axi_wready
	wire          mm_interconnect_0_axi_ad9144_dma_s_axi_awready;                     // axi_ad9144_dma:s_axi_awready -> mm_interconnect_0:axi_ad9144_dma_s_axi_awready
	wire          mm_interconnect_0_axi_ad9144_dma_s_axi_rready;                      // mm_interconnect_0:axi_ad9144_dma_s_axi_rready -> axi_ad9144_dma:s_axi_rready
	wire          mm_interconnect_0_axi_ad9144_dma_s_axi_bready;                      // mm_interconnect_0:axi_ad9144_dma_s_axi_bready -> axi_ad9144_dma:s_axi_bready
	wire          mm_interconnect_0_axi_ad9144_dma_s_axi_wvalid;                      // mm_interconnect_0:axi_ad9144_dma_s_axi_wvalid -> axi_ad9144_dma:s_axi_wvalid
	wire   [11:0] mm_interconnect_0_axi_ad9144_dma_s_axi_araddr;                      // mm_interconnect_0:axi_ad9144_dma_s_axi_araddr -> axi_ad9144_dma:s_axi_araddr
	wire    [2:0] mm_interconnect_0_axi_ad9144_dma_s_axi_arprot;                      // mm_interconnect_0:axi_ad9144_dma_s_axi_arprot -> axi_ad9144_dma:s_axi_arprot
	wire    [1:0] mm_interconnect_0_axi_ad9144_dma_s_axi_rresp;                       // axi_ad9144_dma:s_axi_rresp -> mm_interconnect_0:axi_ad9144_dma_s_axi_rresp
	wire    [2:0] mm_interconnect_0_axi_ad9144_dma_s_axi_awprot;                      // mm_interconnect_0:axi_ad9144_dma_s_axi_awprot -> axi_ad9144_dma:s_axi_awprot
	wire   [31:0] mm_interconnect_0_axi_ad9144_dma_s_axi_wdata;                       // mm_interconnect_0:axi_ad9144_dma_s_axi_wdata -> axi_ad9144_dma:s_axi_wdata
	wire          mm_interconnect_0_axi_ad9144_dma_s_axi_arvalid;                     // mm_interconnect_0:axi_ad9144_dma_s_axi_arvalid -> axi_ad9144_dma:s_axi_arvalid
	wire          mm_interconnect_0_axi_ad9144_dma_s_axi_bvalid;                      // axi_ad9144_dma:s_axi_bvalid -> mm_interconnect_0:axi_ad9144_dma_s_axi_bvalid
	wire          mm_interconnect_0_axi_ad9144_dma_s_axi_awvalid;                     // mm_interconnect_0:axi_ad9144_dma_s_axi_awvalid -> axi_ad9144_dma:s_axi_awvalid
	wire          mm_interconnect_0_axi_ad9144_dma_s_axi_rvalid;                      // axi_ad9144_dma:s_axi_rvalid -> mm_interconnect_0:axi_ad9144_dma_s_axi_rvalid
	wire   [11:0] mm_interconnect_0_axi_ad9680_dma_s_axi_awaddr;                      // mm_interconnect_0:axi_ad9680_dma_s_axi_awaddr -> axi_ad9680_dma:s_axi_awaddr
	wire    [1:0] mm_interconnect_0_axi_ad9680_dma_s_axi_bresp;                       // axi_ad9680_dma:s_axi_bresp -> mm_interconnect_0:axi_ad9680_dma_s_axi_bresp
	wire          mm_interconnect_0_axi_ad9680_dma_s_axi_arready;                     // axi_ad9680_dma:s_axi_arready -> mm_interconnect_0:axi_ad9680_dma_s_axi_arready
	wire   [31:0] mm_interconnect_0_axi_ad9680_dma_s_axi_rdata;                       // axi_ad9680_dma:s_axi_rdata -> mm_interconnect_0:axi_ad9680_dma_s_axi_rdata
	wire    [3:0] mm_interconnect_0_axi_ad9680_dma_s_axi_wstrb;                       // mm_interconnect_0:axi_ad9680_dma_s_axi_wstrb -> axi_ad9680_dma:s_axi_wstrb
	wire          mm_interconnect_0_axi_ad9680_dma_s_axi_wready;                      // axi_ad9680_dma:s_axi_wready -> mm_interconnect_0:axi_ad9680_dma_s_axi_wready
	wire          mm_interconnect_0_axi_ad9680_dma_s_axi_awready;                     // axi_ad9680_dma:s_axi_awready -> mm_interconnect_0:axi_ad9680_dma_s_axi_awready
	wire          mm_interconnect_0_axi_ad9680_dma_s_axi_rready;                      // mm_interconnect_0:axi_ad9680_dma_s_axi_rready -> axi_ad9680_dma:s_axi_rready
	wire          mm_interconnect_0_axi_ad9680_dma_s_axi_bready;                      // mm_interconnect_0:axi_ad9680_dma_s_axi_bready -> axi_ad9680_dma:s_axi_bready
	wire          mm_interconnect_0_axi_ad9680_dma_s_axi_wvalid;                      // mm_interconnect_0:axi_ad9680_dma_s_axi_wvalid -> axi_ad9680_dma:s_axi_wvalid
	wire   [11:0] mm_interconnect_0_axi_ad9680_dma_s_axi_araddr;                      // mm_interconnect_0:axi_ad9680_dma_s_axi_araddr -> axi_ad9680_dma:s_axi_araddr
	wire    [2:0] mm_interconnect_0_axi_ad9680_dma_s_axi_arprot;                      // mm_interconnect_0:axi_ad9680_dma_s_axi_arprot -> axi_ad9680_dma:s_axi_arprot
	wire    [1:0] mm_interconnect_0_axi_ad9680_dma_s_axi_rresp;                       // axi_ad9680_dma:s_axi_rresp -> mm_interconnect_0:axi_ad9680_dma_s_axi_rresp
	wire    [2:0] mm_interconnect_0_axi_ad9680_dma_s_axi_awprot;                      // mm_interconnect_0:axi_ad9680_dma_s_axi_awprot -> axi_ad9680_dma:s_axi_awprot
	wire   [31:0] mm_interconnect_0_axi_ad9680_dma_s_axi_wdata;                       // mm_interconnect_0:axi_ad9680_dma_s_axi_wdata -> axi_ad9680_dma:s_axi_wdata
	wire          mm_interconnect_0_axi_ad9680_dma_s_axi_arvalid;                     // mm_interconnect_0:axi_ad9680_dma_s_axi_arvalid -> axi_ad9680_dma:s_axi_arvalid
	wire          mm_interconnect_0_axi_ad9680_dma_s_axi_bvalid;                      // axi_ad9680_dma:s_axi_bvalid -> mm_interconnect_0:axi_ad9680_dma_s_axi_bvalid
	wire          mm_interconnect_0_axi_ad9680_dma_s_axi_awvalid;                     // mm_interconnect_0:axi_ad9680_dma_s_axi_awvalid -> axi_ad9680_dma:s_axi_awvalid
	wire          mm_interconnect_0_axi_ad9680_dma_s_axi_rvalid;                      // axi_ad9680_dma:s_axi_rvalid -> mm_interconnect_0:axi_ad9680_dma_s_axi_rvalid
	wire          mm_interconnect_0_sys_spi_spi_control_port_chipselect;              // mm_interconnect_0:sys_spi_spi_control_port_chipselect -> sys_spi:spi_select
	wire   [15:0] mm_interconnect_0_sys_spi_spi_control_port_readdata;                // sys_spi:data_to_cpu -> mm_interconnect_0:sys_spi_spi_control_port_readdata
	wire    [2:0] mm_interconnect_0_sys_spi_spi_control_port_address;                 // mm_interconnect_0:sys_spi_spi_control_port_address -> sys_spi:mem_addr
	wire          mm_interconnect_0_sys_spi_spi_control_port_read;                    // mm_interconnect_0:sys_spi_spi_control_port_read -> sys_spi:read_n
	wire          mm_interconnect_0_sys_spi_spi_control_port_write;                   // mm_interconnect_0:sys_spi_spi_control_port_write -> sys_spi:write_n
	wire   [15:0] mm_interconnect_0_sys_spi_spi_control_port_writedata;               // mm_interconnect_0:sys_spi_spi_control_port_writedata -> sys_spi:data_from_cpu
	wire   [31:0] mm_interconnect_0_sys_flash_uas_readdata;                           // sys_flash:uas_readdata -> mm_interconnect_0:sys_flash_uas_readdata
	wire          mm_interconnect_0_sys_flash_uas_waitrequest;                        // sys_flash:uas_waitrequest -> mm_interconnect_0:sys_flash_uas_waitrequest
	wire          mm_interconnect_0_sys_flash_uas_debugaccess;                        // mm_interconnect_0:sys_flash_uas_debugaccess -> sys_flash:uas_debugaccess
	wire   [23:0] mm_interconnect_0_sys_flash_uas_address;                            // mm_interconnect_0:sys_flash_uas_address -> sys_flash:uas_address
	wire          mm_interconnect_0_sys_flash_uas_read;                               // mm_interconnect_0:sys_flash_uas_read -> sys_flash:uas_read
	wire    [3:0] mm_interconnect_0_sys_flash_uas_byteenable;                         // mm_interconnect_0:sys_flash_uas_byteenable -> sys_flash:uas_byteenable
	wire          mm_interconnect_0_sys_flash_uas_readdatavalid;                      // sys_flash:uas_readdatavalid -> mm_interconnect_0:sys_flash_uas_readdatavalid
	wire          mm_interconnect_0_sys_flash_uas_lock;                               // mm_interconnect_0:sys_flash_uas_lock -> sys_flash:uas_lock
	wire          mm_interconnect_0_sys_flash_uas_write;                              // mm_interconnect_0:sys_flash_uas_write -> sys_flash:uas_write
	wire   [31:0] mm_interconnect_0_sys_flash_uas_writedata;                          // mm_interconnect_0:sys_flash_uas_writedata -> sys_flash:uas_writedata
	wire    [2:0] mm_interconnect_0_sys_flash_uas_burstcount;                         // mm_interconnect_0:sys_flash_uas_burstcount -> sys_flash:uas_burstcount
	wire   [31:0] sys_cpu_tightly_coupled_data_master_0_readdata;                     // mm_interconnect_1:sys_cpu_tightly_coupled_data_master_0_readdata -> sys_cpu:dtcm0_readdata
	wire   [28:0] sys_cpu_tightly_coupled_data_master_0_address;                      // sys_cpu:dtcm0_address -> mm_interconnect_1:sys_cpu_tightly_coupled_data_master_0_address
	wire          sys_cpu_tightly_coupled_data_master_0_read;                         // sys_cpu:dtcm0_read -> mm_interconnect_1:sys_cpu_tightly_coupled_data_master_0_read
	wire    [3:0] sys_cpu_tightly_coupled_data_master_0_byteenable;                   // sys_cpu:dtcm0_byteenable -> mm_interconnect_1:sys_cpu_tightly_coupled_data_master_0_byteenable
	wire          sys_cpu_tightly_coupled_data_master_0_write;                        // sys_cpu:dtcm0_write -> mm_interconnect_1:sys_cpu_tightly_coupled_data_master_0_write
	wire   [31:0] sys_cpu_tightly_coupled_data_master_0_writedata;                    // sys_cpu:dtcm0_writedata -> mm_interconnect_1:sys_cpu_tightly_coupled_data_master_0_writedata
	wire          mm_interconnect_1_sys_tlb_mem_s1_chipselect;                        // mm_interconnect_1:sys_tlb_mem_s1_chipselect -> sys_tlb_mem:chipselect
	wire   [31:0] mm_interconnect_1_sys_tlb_mem_s1_readdata;                          // sys_tlb_mem:readdata -> mm_interconnect_1:sys_tlb_mem_s1_readdata
	wire   [15:0] mm_interconnect_1_sys_tlb_mem_s1_address;                           // mm_interconnect_1:sys_tlb_mem_s1_address -> sys_tlb_mem:address
	wire    [3:0] mm_interconnect_1_sys_tlb_mem_s1_byteenable;                        // mm_interconnect_1:sys_tlb_mem_s1_byteenable -> sys_tlb_mem:byteenable
	wire          mm_interconnect_1_sys_tlb_mem_s1_write;                             // mm_interconnect_1:sys_tlb_mem_s1_write -> sys_tlb_mem:write
	wire   [31:0] mm_interconnect_1_sys_tlb_mem_s1_writedata;                         // mm_interconnect_1:sys_tlb_mem_s1_writedata -> sys_tlb_mem:writedata
	wire          mm_interconnect_1_sys_tlb_mem_s1_clken;                             // mm_interconnect_1:sys_tlb_mem_s1_clken -> sys_tlb_mem:clken
	wire   [31:0] sys_cpu_tightly_coupled_instruction_master_0_readdata;              // mm_interconnect_2:sys_cpu_tightly_coupled_instruction_master_0_readdata -> sys_cpu:itcm0_readdata
	wire   [28:0] sys_cpu_tightly_coupled_instruction_master_0_address;               // sys_cpu:itcm0_address -> mm_interconnect_2:sys_cpu_tightly_coupled_instruction_master_0_address
	wire          sys_cpu_tightly_coupled_instruction_master_0_read;                  // sys_cpu:itcm0_read -> mm_interconnect_2:sys_cpu_tightly_coupled_instruction_master_0_read
	wire          mm_interconnect_2_sys_tlb_mem_s2_chipselect;                        // mm_interconnect_2:sys_tlb_mem_s2_chipselect -> sys_tlb_mem:chipselect2
	wire   [31:0] mm_interconnect_2_sys_tlb_mem_s2_readdata;                          // sys_tlb_mem:readdata2 -> mm_interconnect_2:sys_tlb_mem_s2_readdata
	wire   [15:0] mm_interconnect_2_sys_tlb_mem_s2_address;                           // mm_interconnect_2:sys_tlb_mem_s2_address -> sys_tlb_mem:address2
	wire    [3:0] mm_interconnect_2_sys_tlb_mem_s2_byteenable;                        // mm_interconnect_2:sys_tlb_mem_s2_byteenable -> sys_tlb_mem:byteenable2
	wire          mm_interconnect_2_sys_tlb_mem_s2_write;                             // mm_interconnect_2:sys_tlb_mem_s2_write -> sys_tlb_mem:write2
	wire   [31:0] mm_interconnect_2_sys_tlb_mem_s2_writedata;                         // mm_interconnect_2:sys_tlb_mem_s2_writedata -> sys_tlb_mem:writedata2
	wire          mm_interconnect_2_sys_tlb_mem_s2_clken;                             // mm_interconnect_2:sys_tlb_mem_s2_clken -> sys_tlb_mem:clken2
	wire          irq_mapper_receiver0_irq;                                           // sys_ethernet_dma_rx:csr_irq_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                           // sys_ethernet_dma_tx:csr_irq_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                           // axi_ad9680_dma:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                           // axi_ad9144_dma:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                           // sys_uart:av_irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                           // sys_timer_2:irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                           // sys_timer_1:irq -> irq_mapper:receiver6_irq
	wire          irq_mapper_receiver7_irq;                                           // sys_gpio_in:irq -> irq_mapper:receiver7_irq
	wire          irq_mapper_receiver8_irq;                                           // sys_gpio_bd:irq -> irq_mapper:receiver8_irq
	wire          irq_mapper_receiver9_irq;                                           // sys_spi:irq -> irq_mapper:receiver9_irq
	wire   [31:0] sys_cpu_irq_irq;                                                    // irq_mapper:sender_irq -> sys_cpu:irq
	wire          sys_ethernet_receive_valid;                                         // sys_ethernet:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire   [31:0] sys_ethernet_receive_data;                                          // sys_ethernet:ff_rx_data -> avalon_st_adapter:in_0_data
	wire          sys_ethernet_receive_ready;                                         // avalon_st_adapter:in_0_ready -> sys_ethernet:ff_rx_rdy
	wire          sys_ethernet_receive_startofpacket;                                 // sys_ethernet:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire          sys_ethernet_receive_endofpacket;                                   // sys_ethernet:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire    [5:0] sys_ethernet_receive_error;                                         // sys_ethernet:rx_err -> avalon_st_adapter:in_0_error
	wire    [1:0] sys_ethernet_receive_empty;                                         // sys_ethernet:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire          avalon_st_adapter_out_0_valid;                                      // avalon_st_adapter:out_0_valid -> sys_ethernet_dma_rx:st_sink_valid
	wire   [63:0] avalon_st_adapter_out_0_data;                                       // avalon_st_adapter:out_0_data -> sys_ethernet_dma_rx:st_sink_data
	wire          avalon_st_adapter_out_0_ready;                                      // sys_ethernet_dma_rx:st_sink_ready -> avalon_st_adapter:out_0_ready
	wire          avalon_st_adapter_out_0_startofpacket;                              // avalon_st_adapter:out_0_startofpacket -> sys_ethernet_dma_rx:st_sink_startofpacket
	wire          avalon_st_adapter_out_0_endofpacket;                                // avalon_st_adapter:out_0_endofpacket -> sys_ethernet_dma_rx:st_sink_endofpacket
	wire    [5:0] avalon_st_adapter_out_0_error;                                      // avalon_st_adapter:out_0_error -> sys_ethernet_dma_rx:st_sink_error
	wire    [2:0] avalon_st_adapter_out_0_empty;                                      // avalon_st_adapter:out_0_empty -> sys_ethernet_dma_rx:st_sink_empty
	wire          sys_ethernet_dma_tx_st_source_valid;                                // sys_ethernet_dma_tx:st_source_valid -> avalon_st_adapter_001:in_0_valid
	wire   [63:0] sys_ethernet_dma_tx_st_source_data;                                 // sys_ethernet_dma_tx:st_source_data -> avalon_st_adapter_001:in_0_data
	wire          sys_ethernet_dma_tx_st_source_ready;                                // avalon_st_adapter_001:in_0_ready -> sys_ethernet_dma_tx:st_source_ready
	wire          sys_ethernet_dma_tx_st_source_startofpacket;                        // sys_ethernet_dma_tx:st_source_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	wire          sys_ethernet_dma_tx_st_source_endofpacket;                          // sys_ethernet_dma_tx:st_source_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	wire          sys_ethernet_dma_tx_st_source_error;                                // sys_ethernet_dma_tx:st_source_error -> avalon_st_adapter_001:in_0_error
	wire    [2:0] sys_ethernet_dma_tx_st_source_empty;                                // sys_ethernet_dma_tx:st_source_empty -> avalon_st_adapter_001:in_0_empty
	wire          avalon_st_adapter_001_out_0_valid;                                  // avalon_st_adapter_001:out_0_valid -> sys_ethernet:ff_tx_wren
	wire   [31:0] avalon_st_adapter_001_out_0_data;                                   // avalon_st_adapter_001:out_0_data -> sys_ethernet:ff_tx_data
	wire          avalon_st_adapter_001_out_0_ready;                                  // sys_ethernet:ff_tx_rdy -> avalon_st_adapter_001:out_0_ready
	wire          avalon_st_adapter_001_out_0_startofpacket;                          // avalon_st_adapter_001:out_0_startofpacket -> sys_ethernet:ff_tx_sop
	wire          avalon_st_adapter_001_out_0_endofpacket;                            // avalon_st_adapter_001:out_0_endofpacket -> sys_ethernet:ff_tx_eop
	wire          avalon_st_adapter_001_out_0_error;                                  // avalon_st_adapter_001:out_0_error -> sys_ethernet:ff_tx_err
	wire    [1:0] avalon_st_adapter_001_out_0_empty;                                  // avalon_st_adapter_001:out_0_empty -> sys_ethernet:ff_tx_mod
	wire          rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [ad9144_jesd204:sys_resetn_reset_n, ad9680_jesd204:sys_resetn_reset_n, avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, avl_adxcfg_0:rcfg_reset_n, avl_adxcfg_1:rcfg_reset_n, avl_adxcfg_2:rcfg_reset_n, avl_adxcfg_3:rcfg_reset_n, axi_ad9144_dma:s_axi_aresetn, axi_ad9680_dma:s_axi_aresetn, mm_interconnect_0:axi_ad9680_dma_s_axi_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sys_tlb_mem_reset1_reset_bridge_in_reset_reset, mm_interconnect_2:sys_tlb_mem_reset2_reset_bridge_in_reset_reset, rst_translator:in_reset, sys_ethernet:reset, sys_ethernet_reset:in_reset, sys_flash:reset_reset, sys_flash_bridge:reset, sys_gpio_bd:reset_n, sys_gpio_in:reset_n, sys_gpio_out:reset_n, sys_id:reset_n, sys_int_mem:reset, sys_spi:reset_n, sys_timer_1:reset_n, sys_timer_2:reset_n, sys_tlb_mem:reset, sys_tlb_mem:reset2, sys_uart:rst_n]
	wire          rst_controller_reset_out_reset_req;                                 // rst_controller:reset_req -> [rst_translator:reset_req_in, sys_int_mem:reset_req, sys_tlb_mem:reset_req, sys_tlb_mem:reset_req2]
	wire          rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> ad9680_adcfifo:adc_rst
	wire          sys_dma_clk_clk_reset_reset;                                        // sys_dma_clk:reset_n_out -> [rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	wire          rst_controller_002_reset_out_reset;                                 // rst_controller_002:reset_out -> [avl_ad9144_fifo:dma_rst, axi_ad9144_dma:m_src_axi_aresetn, axi_ad9680_dma:m_dest_axi_aresetn, mm_interconnect_0:axi_ad9680_dma_m_dest_axi_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_003_reset_out_reset;                                 // rst_controller_003:reset_out -> avl_ad9144_fifo:dac_rst
	wire          ad9144_jesd204_link_reset_reset;                                    // ad9144_jesd204:link_reset_reset -> rst_controller_003:reset_in0
	wire          rst_controller_004_reset_out_reset;                                 // rst_controller_004:reset_out -> [irq_mapper:reset, mm_interconnect_0:sys_cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sys_cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_2:sys_cpu_reset_reset_bridge_in_reset_reset, rst_translator_001:in_reset, sys_cpu:reset_n]
	wire          rst_controller_004_reset_out_reset_req;                             // rst_controller_004:reset_req -> [rst_translator_001:reset_req_in, sys_cpu:reset_req]
	wire          sys_cpu_debug_reset_request_reset;                                  // sys_cpu:debug_reset_request -> rst_controller_004:reset_in1
	wire          rst_controller_005_reset_out_reset;                                 // rst_controller_005:reset_out -> [sys_ethernet_dma_rx:reset_n_reset_n, sys_ethernet_dma_tx:reset_n_reset_n]
	wire          rst_controller_006_reset_out_reset;                                 // rst_controller_006:reset_out -> mm_interconnect_0:sys_ddr3_cntrl_ctrl_amm_0_translator_reset_reset_bridge_in_reset_reset

	system_bd_ad9144_jesd204 ad9144_jesd204 (
		.sys_clk_clk        (sys_clk_clk_clk),                 //   input,  width = 1,    sys_clk.clk
		.sys_resetn_reset_n (~rst_controller_reset_out_reset), //   input,  width = 1, sys_resetn.reset_n
		.ref_clk_clk        (tx_ref_clk_clk),                  //   input,  width = 1,    ref_clk.clk
		.link_clk_clk       (ad9144_jesd204_link_clk_clk),     //  output,  width = 1,   link_clk.clk
		.link_reset_reset   (ad9144_jesd204_link_reset_reset)  //  output,  width = 1, link_reset.reset
	);

	system_bd_ad9680_adcfifo ad9680_adcfifo (
		.adc_clk         (ad9680_jesd204_link_clk_clk),                //   input,    width = 1,         if_adc_clk.clk
		.adc_rst         (rst_controller_001_reset_out_reset),         //   input,    width = 1,         if_adc_rst.reset
		.adc_wr          (),                                           //   input,    width = 1,          if_adc_wr.valid
		.adc_wdata       (),                                           //   input,  width = 128,       if_adc_wdata.data
		.adc_wovf        (),                                           //  output,    width = 1,        if_adc_wovf.ovf
		.dma_clk         (sys_dma_clk_clk_clk),                        //   input,    width = 1,         if_dma_clk.clk
		.dma_wr          (ad9680_adcfifo_if_dma_wr_valid),             //  output,    width = 1,          if_dma_wr.valid
		.dma_wdata       (ad9680_adcfifo_if_dma_wdata_data),           //  output,  width = 128,       if_dma_wdata.data
		.dma_wready      (axi_ad9680_dma_if_s_axis_ready_ready),       //   input,    width = 1,      if_dma_wready.ready
		.dma_xfer_req    (axi_ad9680_dma_if_s_axis_xfer_req_xfer_req), //   input,    width = 1,    if_dma_xfer_req.xfer_req
		.dma_xfer_status ()                                            //  output,    width = 4, if_dma_xfer_status.xfer_status
	);

	system_bd_ad9680_jesd204 ad9680_jesd204 (
		.sys_clk_clk        (sys_clk_clk_clk),                 //   input,  width = 1,    sys_clk.clk
		.sys_resetn_reset_n (~rst_controller_reset_out_reset), //   input,  width = 1, sys_resetn.reset_n
		.ref_clk_clk        (rx_ref_clk_clk),                  //   input,  width = 1,    ref_clk.clk
		.link_clk_clk       (ad9680_jesd204_link_clk_clk),     //  output,  width = 1,   link_clk.clk
		.link_reset_reset   ()                                 //  output,  width = 1, link_reset.reset
	);

	system_bd_avl_ad9144_fifo avl_ad9144_fifo (
		.dma_clk       (sys_dma_clk_clk_clk),                        //   input,    width = 1,       if_dma_clk.clk
		.dma_rst       (rst_controller_002_reset_out_reset),         //   input,    width = 1,       if_dma_rst.reset
		.dma_valid     (axi_ad9144_dma_if_m_axis_valid_valid),       //   input,    width = 1,     if_dma_valid.valid
		.dma_data      (axi_ad9144_dma_if_m_axis_data_data),         //   input,  width = 128,      if_dma_data.data
		.dma_ready     (avl_ad9144_fifo_if_dma_ready_ready),         //  output,    width = 1,     if_dma_ready.ready
		.dma_xfer_req  (axi_ad9144_dma_if_m_axis_xfer_req_xfer_req), //   input,    width = 1,  if_dma_xfer_req.xfer_req
		.dma_xfer_last (axi_ad9144_dma_if_m_axis_last_last),         //   input,    width = 1, if_dma_xfer_last.last
		.dac_clk       (ad9144_jesd204_link_clk_clk),                //   input,    width = 1,       if_dac_clk.clk
		.dac_rst       (rst_controller_003_reset_out_reset),         //   input,    width = 1,       if_dac_rst.reset
		.dac_valid     (util_ad9144_upack_if_dac_valid_valid),       //   input,    width = 1,     if_dac_valid.valid
		.dac_data      (avl_ad9144_fifo_if_dac_data_data),           //  output,  width = 128,      if_dac_data.data
		.dac_xfer_out  (),                                           //  output,    width = 1,  if_dac_xfer_out.xfer_req
		.dac_dunf      (),                                           //  output,    width = 1,      if_dac_dunf.unf
		.bypass        (tx_fifo_bypass_bypass)                       //   input,    width = 1,        if_bypass.bypass
	);

	system_bd_avl_adxcfg_0 avl_adxcfg_0 (
		.rcfg_clk               (sys_clk_clk_clk),                                    //   input,   width = 1,     rcfg_clk.clk
		.rcfg_reset_n           (~rst_controller_reset_out_reset),                    //   input,   width = 1, rcfg_reset_n.reset_n
		.rcfg_in_read_0         (mm_interconnect_0_avl_adxcfg_0_rcfg_s0_read),        //   input,   width = 1,      rcfg_s0.read
		.rcfg_in_write_0        (mm_interconnect_0_avl_adxcfg_0_rcfg_s0_write),       //   input,   width = 1,             .write
		.rcfg_in_address_0      (mm_interconnect_0_avl_adxcfg_0_rcfg_s0_address),     //   input,  width = 10,             .address
		.rcfg_in_writedata_0    (mm_interconnect_0_avl_adxcfg_0_rcfg_s0_writedata),   //   input,  width = 32,             .writedata
		.rcfg_in_readdata_0     (mm_interconnect_0_avl_adxcfg_0_rcfg_s0_readdata),    //  output,  width = 32,             .readdata
		.rcfg_in_waitrequest_0  (mm_interconnect_0_avl_adxcfg_0_rcfg_s0_waitrequest), //  output,   width = 1,             .waitrequest
		.rcfg_out_read_0        (),                                                   //  output,   width = 1,      rcfg_m0.read
		.rcfg_out_write_0       (),                                                   //  output,   width = 1,             .write
		.rcfg_out_address_0     (),                                                   //  output,  width = 10,             .address
		.rcfg_out_writedata_0   (),                                                   //  output,  width = 32,             .writedata
		.rcfg_out_readdata_0    (),                                                   //   input,  width = 32,             .readdata
		.rcfg_out_waitrequest_0 (),                                                   //   input,   width = 1,             .waitrequest
		.rcfg_in_read_1         (mm_interconnect_0_avl_adxcfg_0_rcfg_s1_read),        //   input,   width = 1,      rcfg_s1.read
		.rcfg_in_write_1        (mm_interconnect_0_avl_adxcfg_0_rcfg_s1_write),       //   input,   width = 1,             .write
		.rcfg_in_address_1      (mm_interconnect_0_avl_adxcfg_0_rcfg_s1_address),     //   input,  width = 10,             .address
		.rcfg_in_writedata_1    (mm_interconnect_0_avl_adxcfg_0_rcfg_s1_writedata),   //   input,  width = 32,             .writedata
		.rcfg_in_readdata_1     (mm_interconnect_0_avl_adxcfg_0_rcfg_s1_readdata),    //  output,  width = 32,             .readdata
		.rcfg_in_waitrequest_1  (mm_interconnect_0_avl_adxcfg_0_rcfg_s1_waitrequest), //  output,   width = 1,             .waitrequest
		.rcfg_out_read_1        (),                                                   //  output,   width = 1,      rcfg_m1.read
		.rcfg_out_write_1       (),                                                   //  output,   width = 1,             .write
		.rcfg_out_address_1     (),                                                   //  output,  width = 10,             .address
		.rcfg_out_writedata_1   (),                                                   //  output,  width = 32,             .writedata
		.rcfg_out_readdata_1    (),                                                   //   input,  width = 32,             .readdata
		.rcfg_out_waitrequest_1 ()                                                    //   input,   width = 1,             .waitrequest
	);

	system_bd_avl_adxcfg_1 avl_adxcfg_1 (
		.rcfg_clk               (sys_clk_clk_clk),                                    //   input,   width = 1,     rcfg_clk.clk
		.rcfg_reset_n           (~rst_controller_reset_out_reset),                    //   input,   width = 1, rcfg_reset_n.reset_n
		.rcfg_in_read_0         (mm_interconnect_0_avl_adxcfg_1_rcfg_s0_read),        //   input,   width = 1,      rcfg_s0.read
		.rcfg_in_write_0        (mm_interconnect_0_avl_adxcfg_1_rcfg_s0_write),       //   input,   width = 1,             .write
		.rcfg_in_address_0      (mm_interconnect_0_avl_adxcfg_1_rcfg_s0_address),     //   input,  width = 10,             .address
		.rcfg_in_writedata_0    (mm_interconnect_0_avl_adxcfg_1_rcfg_s0_writedata),   //   input,  width = 32,             .writedata
		.rcfg_in_readdata_0     (mm_interconnect_0_avl_adxcfg_1_rcfg_s0_readdata),    //  output,  width = 32,             .readdata
		.rcfg_in_waitrequest_0  (mm_interconnect_0_avl_adxcfg_1_rcfg_s0_waitrequest), //  output,   width = 1,             .waitrequest
		.rcfg_out_read_0        (),                                                   //  output,   width = 1,      rcfg_m0.read
		.rcfg_out_write_0       (),                                                   //  output,   width = 1,             .write
		.rcfg_out_address_0     (),                                                   //  output,  width = 10,             .address
		.rcfg_out_writedata_0   (),                                                   //  output,  width = 32,             .writedata
		.rcfg_out_readdata_0    (),                                                   //   input,  width = 32,             .readdata
		.rcfg_out_waitrequest_0 (),                                                   //   input,   width = 1,             .waitrequest
		.rcfg_in_read_1         (mm_interconnect_0_avl_adxcfg_1_rcfg_s1_read),        //   input,   width = 1,      rcfg_s1.read
		.rcfg_in_write_1        (mm_interconnect_0_avl_adxcfg_1_rcfg_s1_write),       //   input,   width = 1,             .write
		.rcfg_in_address_1      (mm_interconnect_0_avl_adxcfg_1_rcfg_s1_address),     //   input,  width = 10,             .address
		.rcfg_in_writedata_1    (mm_interconnect_0_avl_adxcfg_1_rcfg_s1_writedata),   //   input,  width = 32,             .writedata
		.rcfg_in_readdata_1     (mm_interconnect_0_avl_adxcfg_1_rcfg_s1_readdata),    //  output,  width = 32,             .readdata
		.rcfg_in_waitrequest_1  (mm_interconnect_0_avl_adxcfg_1_rcfg_s1_waitrequest), //  output,   width = 1,             .waitrequest
		.rcfg_out_read_1        (),                                                   //  output,   width = 1,      rcfg_m1.read
		.rcfg_out_write_1       (),                                                   //  output,   width = 1,             .write
		.rcfg_out_address_1     (),                                                   //  output,  width = 10,             .address
		.rcfg_out_writedata_1   (),                                                   //  output,  width = 32,             .writedata
		.rcfg_out_readdata_1    (),                                                   //   input,  width = 32,             .readdata
		.rcfg_out_waitrequest_1 ()                                                    //   input,   width = 1,             .waitrequest
	);

	system_bd_avl_adxcfg_2 avl_adxcfg_2 (
		.rcfg_clk               (sys_clk_clk_clk),                                    //   input,   width = 1,     rcfg_clk.clk
		.rcfg_reset_n           (~rst_controller_reset_out_reset),                    //   input,   width = 1, rcfg_reset_n.reset_n
		.rcfg_in_read_0         (mm_interconnect_0_avl_adxcfg_2_rcfg_s0_read),        //   input,   width = 1,      rcfg_s0.read
		.rcfg_in_write_0        (mm_interconnect_0_avl_adxcfg_2_rcfg_s0_write),       //   input,   width = 1,             .write
		.rcfg_in_address_0      (mm_interconnect_0_avl_adxcfg_2_rcfg_s0_address),     //   input,  width = 10,             .address
		.rcfg_in_writedata_0    (mm_interconnect_0_avl_adxcfg_2_rcfg_s0_writedata),   //   input,  width = 32,             .writedata
		.rcfg_in_readdata_0     (mm_interconnect_0_avl_adxcfg_2_rcfg_s0_readdata),    //  output,  width = 32,             .readdata
		.rcfg_in_waitrequest_0  (mm_interconnect_0_avl_adxcfg_2_rcfg_s0_waitrequest), //  output,   width = 1,             .waitrequest
		.rcfg_out_read_0        (),                                                   //  output,   width = 1,      rcfg_m0.read
		.rcfg_out_write_0       (),                                                   //  output,   width = 1,             .write
		.rcfg_out_address_0     (),                                                   //  output,  width = 10,             .address
		.rcfg_out_writedata_0   (),                                                   //  output,  width = 32,             .writedata
		.rcfg_out_readdata_0    (),                                                   //   input,  width = 32,             .readdata
		.rcfg_out_waitrequest_0 (),                                                   //   input,   width = 1,             .waitrequest
		.rcfg_in_read_1         (mm_interconnect_0_avl_adxcfg_2_rcfg_s1_read),        //   input,   width = 1,      rcfg_s1.read
		.rcfg_in_write_1        (mm_interconnect_0_avl_adxcfg_2_rcfg_s1_write),       //   input,   width = 1,             .write
		.rcfg_in_address_1      (mm_interconnect_0_avl_adxcfg_2_rcfg_s1_address),     //   input,  width = 10,             .address
		.rcfg_in_writedata_1    (mm_interconnect_0_avl_adxcfg_2_rcfg_s1_writedata),   //   input,  width = 32,             .writedata
		.rcfg_in_readdata_1     (mm_interconnect_0_avl_adxcfg_2_rcfg_s1_readdata),    //  output,  width = 32,             .readdata
		.rcfg_in_waitrequest_1  (mm_interconnect_0_avl_adxcfg_2_rcfg_s1_waitrequest), //  output,   width = 1,             .waitrequest
		.rcfg_out_read_1        (),                                                   //  output,   width = 1,      rcfg_m1.read
		.rcfg_out_write_1       (),                                                   //  output,   width = 1,             .write
		.rcfg_out_address_1     (),                                                   //  output,  width = 10,             .address
		.rcfg_out_writedata_1   (),                                                   //  output,  width = 32,             .writedata
		.rcfg_out_readdata_1    (),                                                   //   input,  width = 32,             .readdata
		.rcfg_out_waitrequest_1 ()                                                    //   input,   width = 1,             .waitrequest
	);

	system_bd_avl_adxcfg_3 avl_adxcfg_3 (
		.rcfg_clk               (sys_clk_clk_clk),                                    //   input,   width = 1,     rcfg_clk.clk
		.rcfg_reset_n           (~rst_controller_reset_out_reset),                    //   input,   width = 1, rcfg_reset_n.reset_n
		.rcfg_in_read_0         (mm_interconnect_0_avl_adxcfg_3_rcfg_s0_read),        //   input,   width = 1,      rcfg_s0.read
		.rcfg_in_write_0        (mm_interconnect_0_avl_adxcfg_3_rcfg_s0_write),       //   input,   width = 1,             .write
		.rcfg_in_address_0      (mm_interconnect_0_avl_adxcfg_3_rcfg_s0_address),     //   input,  width = 10,             .address
		.rcfg_in_writedata_0    (mm_interconnect_0_avl_adxcfg_3_rcfg_s0_writedata),   //   input,  width = 32,             .writedata
		.rcfg_in_readdata_0     (mm_interconnect_0_avl_adxcfg_3_rcfg_s0_readdata),    //  output,  width = 32,             .readdata
		.rcfg_in_waitrequest_0  (mm_interconnect_0_avl_adxcfg_3_rcfg_s0_waitrequest), //  output,   width = 1,             .waitrequest
		.rcfg_out_read_0        (),                                                   //  output,   width = 1,      rcfg_m0.read
		.rcfg_out_write_0       (),                                                   //  output,   width = 1,             .write
		.rcfg_out_address_0     (),                                                   //  output,  width = 10,             .address
		.rcfg_out_writedata_0   (),                                                   //  output,  width = 32,             .writedata
		.rcfg_out_readdata_0    (),                                                   //   input,  width = 32,             .readdata
		.rcfg_out_waitrequest_0 (),                                                   //   input,   width = 1,             .waitrequest
		.rcfg_in_read_1         (mm_interconnect_0_avl_adxcfg_3_rcfg_s1_read),        //   input,   width = 1,      rcfg_s1.read
		.rcfg_in_write_1        (mm_interconnect_0_avl_adxcfg_3_rcfg_s1_write),       //   input,   width = 1,             .write
		.rcfg_in_address_1      (mm_interconnect_0_avl_adxcfg_3_rcfg_s1_address),     //   input,  width = 10,             .address
		.rcfg_in_writedata_1    (mm_interconnect_0_avl_adxcfg_3_rcfg_s1_writedata),   //   input,  width = 32,             .writedata
		.rcfg_in_readdata_1     (mm_interconnect_0_avl_adxcfg_3_rcfg_s1_readdata),    //  output,  width = 32,             .readdata
		.rcfg_in_waitrequest_1  (mm_interconnect_0_avl_adxcfg_3_rcfg_s1_waitrequest), //  output,   width = 1,             .waitrequest
		.rcfg_out_read_1        (),                                                   //  output,   width = 1,      rcfg_m1.read
		.rcfg_out_write_1       (),                                                   //  output,   width = 1,             .write
		.rcfg_out_address_1     (),                                                   //  output,  width = 10,             .address
		.rcfg_out_writedata_1   (),                                                   //  output,  width = 32,             .writedata
		.rcfg_out_readdata_1    (),                                                   //   input,  width = 32,             .readdata
		.rcfg_out_waitrequest_1 ()                                                    //   input,   width = 1,             .waitrequest
	);

	system_bd_axi_ad9144_core axi_ad9144_core (
	);

	system_bd_axi_ad9144_dma axi_ad9144_dma (
		.s_axi_aclk        (sys_clk_clk_clk),                                //   input,    width = 1,        s_axi_clock.clk
		.s_axi_aresetn     (~rst_controller_reset_out_reset),                //   input,    width = 1,        s_axi_reset.reset_n
		.s_axi_awvalid     (mm_interconnect_0_axi_ad9144_dma_s_axi_awvalid), //   input,    width = 1,              s_axi.awvalid
		.s_axi_awaddr      (mm_interconnect_0_axi_ad9144_dma_s_axi_awaddr),  //   input,   width = 12,                   .awaddr
		.s_axi_awprot      (mm_interconnect_0_axi_ad9144_dma_s_axi_awprot),  //   input,    width = 3,                   .awprot
		.s_axi_awready     (mm_interconnect_0_axi_ad9144_dma_s_axi_awready), //  output,    width = 1,                   .awready
		.s_axi_wvalid      (mm_interconnect_0_axi_ad9144_dma_s_axi_wvalid),  //   input,    width = 1,                   .wvalid
		.s_axi_wdata       (mm_interconnect_0_axi_ad9144_dma_s_axi_wdata),   //   input,   width = 32,                   .wdata
		.s_axi_wstrb       (mm_interconnect_0_axi_ad9144_dma_s_axi_wstrb),   //   input,    width = 4,                   .wstrb
		.s_axi_wready      (mm_interconnect_0_axi_ad9144_dma_s_axi_wready),  //  output,    width = 1,                   .wready
		.s_axi_bvalid      (mm_interconnect_0_axi_ad9144_dma_s_axi_bvalid),  //  output,    width = 1,                   .bvalid
		.s_axi_bresp       (mm_interconnect_0_axi_ad9144_dma_s_axi_bresp),   //  output,    width = 2,                   .bresp
		.s_axi_bready      (mm_interconnect_0_axi_ad9144_dma_s_axi_bready),  //   input,    width = 1,                   .bready
		.s_axi_arvalid     (mm_interconnect_0_axi_ad9144_dma_s_axi_arvalid), //   input,    width = 1,                   .arvalid
		.s_axi_araddr      (mm_interconnect_0_axi_ad9144_dma_s_axi_araddr),  //   input,   width = 12,                   .araddr
		.s_axi_arprot      (mm_interconnect_0_axi_ad9144_dma_s_axi_arprot),  //   input,    width = 3,                   .arprot
		.s_axi_arready     (mm_interconnect_0_axi_ad9144_dma_s_axi_arready), //  output,    width = 1,                   .arready
		.s_axi_rvalid      (mm_interconnect_0_axi_ad9144_dma_s_axi_rvalid),  //  output,    width = 1,                   .rvalid
		.s_axi_rresp       (mm_interconnect_0_axi_ad9144_dma_s_axi_rresp),   //  output,    width = 2,                   .rresp
		.s_axi_rdata       (mm_interconnect_0_axi_ad9144_dma_s_axi_rdata),   //  output,   width = 32,                   .rdata
		.s_axi_rready      (mm_interconnect_0_axi_ad9144_dma_s_axi_rready),  //   input,    width = 1,                   .rready
		.irq               (irq_mapper_receiver3_irq),                       //  output,    width = 1,   interrupt_sender.irq
		.m_src_axi_aclk    (sys_dma_clk_clk_clk),                            //   input,    width = 1,    m_src_axi_clock.clk
		.m_src_axi_aresetn (~rst_controller_002_reset_out_reset),            //   input,    width = 1,    m_src_axi_reset.reset_n
		.m_axis_aclk       (sys_dma_clk_clk_clk),                            //   input,    width = 1,     if_m_axis_aclk.clk
		.m_axis_valid      (axi_ad9144_dma_if_m_axis_valid_valid),           //  output,    width = 1,    if_m_axis_valid.valid
		.m_axis_data       (axi_ad9144_dma_if_m_axis_data_data),             //  output,  width = 128,     if_m_axis_data.data
		.m_axis_ready      (avl_ad9144_fifo_if_dma_ready_ready),             //   input,    width = 1,    if_m_axis_ready.ready
		.m_axis_last       (axi_ad9144_dma_if_m_axis_last_last),             //  output,    width = 1,     if_m_axis_last.last
		.m_axis_xfer_req   (axi_ad9144_dma_if_m_axis_xfer_req_xfer_req),     //  output,    width = 1, if_m_axis_xfer_req.xfer_req
		.m_src_axi_awvalid (axi_ad9144_dma_m_src_axi_awvalid),               //  output,    width = 1,          m_src_axi.awvalid
		.m_src_axi_awaddr  (axi_ad9144_dma_m_src_axi_awaddr),                //  output,   width = 32,                   .awaddr
		.m_src_axi_awready (axi_ad9144_dma_m_src_axi_awready),               //   input,    width = 1,                   .awready
		.m_src_axi_wvalid  (axi_ad9144_dma_m_src_axi_wvalid),                //  output,    width = 1,                   .wvalid
		.m_src_axi_wdata   (axi_ad9144_dma_m_src_axi_wdata),                 //  output,  width = 128,                   .wdata
		.m_src_axi_wstrb   (axi_ad9144_dma_m_src_axi_wstrb),                 //  output,   width = 16,                   .wstrb
		.m_src_axi_wready  (axi_ad9144_dma_m_src_axi_wready),                //   input,    width = 1,                   .wready
		.m_src_axi_bvalid  (axi_ad9144_dma_m_src_axi_bvalid),                //   input,    width = 1,                   .bvalid
		.m_src_axi_bresp   (axi_ad9144_dma_m_src_axi_bresp),                 //   input,    width = 2,                   .bresp
		.m_src_axi_bready  (axi_ad9144_dma_m_src_axi_bready),                //  output,    width = 1,                   .bready
		.m_src_axi_arvalid (axi_ad9144_dma_m_src_axi_arvalid),               //  output,    width = 1,                   .arvalid
		.m_src_axi_araddr  (axi_ad9144_dma_m_src_axi_araddr),                //  output,   width = 32,                   .araddr
		.m_src_axi_arready (axi_ad9144_dma_m_src_axi_arready),               //   input,    width = 1,                   .arready
		.m_src_axi_rvalid  (axi_ad9144_dma_m_src_axi_rvalid),                //   input,    width = 1,                   .rvalid
		.m_src_axi_rresp   (axi_ad9144_dma_m_src_axi_rresp),                 //   input,    width = 2,                   .rresp
		.m_src_axi_rdata   (axi_ad9144_dma_m_src_axi_rdata),                 //   input,  width = 128,                   .rdata
		.m_src_axi_rready  (axi_ad9144_dma_m_src_axi_rready),                //  output,    width = 1,                   .rready
		.m_src_axi_awlen   (axi_ad9144_dma_m_src_axi_awlen),                 //  output,    width = 4,                   .awlen
		.m_src_axi_awsize  (axi_ad9144_dma_m_src_axi_awsize),                //  output,    width = 3,                   .awsize
		.m_src_axi_awburst (axi_ad9144_dma_m_src_axi_awburst),               //  output,    width = 2,                   .awburst
		.m_src_axi_awcache (axi_ad9144_dma_m_src_axi_awcache),               //  output,    width = 4,                   .awcache
		.m_src_axi_awprot  (axi_ad9144_dma_m_src_axi_awprot),                //  output,    width = 3,                   .awprot
		.m_src_axi_wlast   (axi_ad9144_dma_m_src_axi_wlast),                 //  output,    width = 1,                   .wlast
		.m_src_axi_arlen   (axi_ad9144_dma_m_src_axi_arlen),                 //  output,    width = 4,                   .arlen
		.m_src_axi_arsize  (axi_ad9144_dma_m_src_axi_arsize),                //  output,    width = 3,                   .arsize
		.m_src_axi_arburst (axi_ad9144_dma_m_src_axi_arburst),               //  output,    width = 2,                   .arburst
		.m_src_axi_arcache (axi_ad9144_dma_m_src_axi_arcache),               //  output,    width = 4,                   .arcache
		.m_src_axi_arprot  (axi_ad9144_dma_m_src_axi_arprot),                //  output,    width = 3,                   .arprot
		.m_src_axi_awid    (axi_ad9144_dma_m_src_axi_awid),                  //  output,    width = 1,                   .awid
		.m_src_axi_awlock  (axi_ad9144_dma_m_src_axi_awlock),                //  output,    width = 2,                   .awlock
		.m_src_axi_wid     (axi_ad9144_dma_m_src_axi_wid),                   //  output,    width = 1,                   .wid
		.m_src_axi_arid    (axi_ad9144_dma_m_src_axi_arid),                  //  output,    width = 1,                   .arid
		.m_src_axi_arlock  (axi_ad9144_dma_m_src_axi_arlock),                //  output,    width = 2,                   .arlock
		.m_src_axi_rid     (axi_ad9144_dma_m_src_axi_rid),                   //   input,    width = 1,                   .rid
		.m_src_axi_bid     (axi_ad9144_dma_m_src_axi_bid),                   //   input,    width = 1,                   .bid
		.m_src_axi_rlast   (axi_ad9144_dma_m_src_axi_rlast)                  //   input,    width = 1,                   .rlast
	);

	system_bd_axi_ad9680_core axi_ad9680_core (
	);

	system_bd_axi_ad9680_dma axi_ad9680_dma (
		.s_axi_aclk         (sys_clk_clk_clk),                                //   input,    width = 1,        s_axi_clock.clk
		.s_axi_aresetn      (~rst_controller_reset_out_reset),                //   input,    width = 1,        s_axi_reset.reset_n
		.s_axi_awvalid      (mm_interconnect_0_axi_ad9680_dma_s_axi_awvalid), //   input,    width = 1,              s_axi.awvalid
		.s_axi_awaddr       (mm_interconnect_0_axi_ad9680_dma_s_axi_awaddr),  //   input,   width = 12,                   .awaddr
		.s_axi_awprot       (mm_interconnect_0_axi_ad9680_dma_s_axi_awprot),  //   input,    width = 3,                   .awprot
		.s_axi_awready      (mm_interconnect_0_axi_ad9680_dma_s_axi_awready), //  output,    width = 1,                   .awready
		.s_axi_wvalid       (mm_interconnect_0_axi_ad9680_dma_s_axi_wvalid),  //   input,    width = 1,                   .wvalid
		.s_axi_wdata        (mm_interconnect_0_axi_ad9680_dma_s_axi_wdata),   //   input,   width = 32,                   .wdata
		.s_axi_wstrb        (mm_interconnect_0_axi_ad9680_dma_s_axi_wstrb),   //   input,    width = 4,                   .wstrb
		.s_axi_wready       (mm_interconnect_0_axi_ad9680_dma_s_axi_wready),  //  output,    width = 1,                   .wready
		.s_axi_bvalid       (mm_interconnect_0_axi_ad9680_dma_s_axi_bvalid),  //  output,    width = 1,                   .bvalid
		.s_axi_bresp        (mm_interconnect_0_axi_ad9680_dma_s_axi_bresp),   //  output,    width = 2,                   .bresp
		.s_axi_bready       (mm_interconnect_0_axi_ad9680_dma_s_axi_bready),  //   input,    width = 1,                   .bready
		.s_axi_arvalid      (mm_interconnect_0_axi_ad9680_dma_s_axi_arvalid), //   input,    width = 1,                   .arvalid
		.s_axi_araddr       (mm_interconnect_0_axi_ad9680_dma_s_axi_araddr),  //   input,   width = 12,                   .araddr
		.s_axi_arprot       (mm_interconnect_0_axi_ad9680_dma_s_axi_arprot),  //   input,    width = 3,                   .arprot
		.s_axi_arready      (mm_interconnect_0_axi_ad9680_dma_s_axi_arready), //  output,    width = 1,                   .arready
		.s_axi_rvalid       (mm_interconnect_0_axi_ad9680_dma_s_axi_rvalid),  //  output,    width = 1,                   .rvalid
		.s_axi_rresp        (mm_interconnect_0_axi_ad9680_dma_s_axi_rresp),   //  output,    width = 2,                   .rresp
		.s_axi_rdata        (mm_interconnect_0_axi_ad9680_dma_s_axi_rdata),   //  output,   width = 32,                   .rdata
		.s_axi_rready       (mm_interconnect_0_axi_ad9680_dma_s_axi_rready),  //   input,    width = 1,                   .rready
		.irq                (irq_mapper_receiver2_irq),                       //  output,    width = 1,   interrupt_sender.irq
		.m_dest_axi_aclk    (sys_dma_clk_clk_clk),                            //   input,    width = 1,   m_dest_axi_clock.clk
		.m_dest_axi_aresetn (~rst_controller_002_reset_out_reset),            //   input,    width = 1,   m_dest_axi_reset.reset_n
		.s_axis_aclk        (sys_dma_clk_clk_clk),                            //   input,    width = 1,     if_s_axis_aclk.clk
		.s_axis_valid       (ad9680_adcfifo_if_dma_wr_valid),                 //   input,    width = 1,    if_s_axis_valid.valid
		.s_axis_data        (ad9680_adcfifo_if_dma_wdata_data),               //   input,  width = 128,     if_s_axis_data.data
		.s_axis_ready       (axi_ad9680_dma_if_s_axis_ready_ready),           //  output,    width = 1,    if_s_axis_ready.ready
		.s_axis_xfer_req    (axi_ad9680_dma_if_s_axis_xfer_req_xfer_req),     //  output,    width = 1, if_s_axis_xfer_req.xfer_req
		.m_dest_axi_awvalid (axi_ad9680_dma_m_dest_axi_awvalid),              //  output,    width = 1,         m_dest_axi.awvalid
		.m_dest_axi_awaddr  (axi_ad9680_dma_m_dest_axi_awaddr),               //  output,   width = 32,                   .awaddr
		.m_dest_axi_awready (axi_ad9680_dma_m_dest_axi_awready),              //   input,    width = 1,                   .awready
		.m_dest_axi_wvalid  (axi_ad9680_dma_m_dest_axi_wvalid),               //  output,    width = 1,                   .wvalid
		.m_dest_axi_wdata   (axi_ad9680_dma_m_dest_axi_wdata),                //  output,  width = 128,                   .wdata
		.m_dest_axi_wstrb   (axi_ad9680_dma_m_dest_axi_wstrb),                //  output,   width = 16,                   .wstrb
		.m_dest_axi_wready  (axi_ad9680_dma_m_dest_axi_wready),               //   input,    width = 1,                   .wready
		.m_dest_axi_bvalid  (axi_ad9680_dma_m_dest_axi_bvalid),               //   input,    width = 1,                   .bvalid
		.m_dest_axi_bresp   (axi_ad9680_dma_m_dest_axi_bresp),                //   input,    width = 2,                   .bresp
		.m_dest_axi_bready  (axi_ad9680_dma_m_dest_axi_bready),               //  output,    width = 1,                   .bready
		.m_dest_axi_arvalid (axi_ad9680_dma_m_dest_axi_arvalid),              //  output,    width = 1,                   .arvalid
		.m_dest_axi_araddr  (axi_ad9680_dma_m_dest_axi_araddr),               //  output,   width = 32,                   .araddr
		.m_dest_axi_arready (axi_ad9680_dma_m_dest_axi_arready),              //   input,    width = 1,                   .arready
		.m_dest_axi_rvalid  (axi_ad9680_dma_m_dest_axi_rvalid),               //   input,    width = 1,                   .rvalid
		.m_dest_axi_rresp   (axi_ad9680_dma_m_dest_axi_rresp),                //   input,    width = 2,                   .rresp
		.m_dest_axi_rdata   (axi_ad9680_dma_m_dest_axi_rdata),                //   input,  width = 128,                   .rdata
		.m_dest_axi_rready  (axi_ad9680_dma_m_dest_axi_rready),               //  output,    width = 1,                   .rready
		.m_dest_axi_awlen   (axi_ad9680_dma_m_dest_axi_awlen),                //  output,    width = 4,                   .awlen
		.m_dest_axi_awsize  (axi_ad9680_dma_m_dest_axi_awsize),               //  output,    width = 3,                   .awsize
		.m_dest_axi_awburst (axi_ad9680_dma_m_dest_axi_awburst),              //  output,    width = 2,                   .awburst
		.m_dest_axi_awcache (axi_ad9680_dma_m_dest_axi_awcache),              //  output,    width = 4,                   .awcache
		.m_dest_axi_awprot  (axi_ad9680_dma_m_dest_axi_awprot),               //  output,    width = 3,                   .awprot
		.m_dest_axi_wlast   (axi_ad9680_dma_m_dest_axi_wlast),                //  output,    width = 1,                   .wlast
		.m_dest_axi_arlen   (axi_ad9680_dma_m_dest_axi_arlen),                //  output,    width = 4,                   .arlen
		.m_dest_axi_arsize  (axi_ad9680_dma_m_dest_axi_arsize),               //  output,    width = 3,                   .arsize
		.m_dest_axi_arburst (axi_ad9680_dma_m_dest_axi_arburst),              //  output,    width = 2,                   .arburst
		.m_dest_axi_arcache (axi_ad9680_dma_m_dest_axi_arcache),              //  output,    width = 4,                   .arcache
		.m_dest_axi_arprot  (axi_ad9680_dma_m_dest_axi_arprot),               //  output,    width = 3,                   .arprot
		.m_dest_axi_awid    (axi_ad9680_dma_m_dest_axi_awid),                 //  output,    width = 1,                   .awid
		.m_dest_axi_awlock  (axi_ad9680_dma_m_dest_axi_awlock),               //  output,    width = 2,                   .awlock
		.m_dest_axi_wid     (axi_ad9680_dma_m_dest_axi_wid),                  //  output,    width = 1,                   .wid
		.m_dest_axi_arid    (axi_ad9680_dma_m_dest_axi_arid),                 //  output,    width = 1,                   .arid
		.m_dest_axi_arlock  (axi_ad9680_dma_m_dest_axi_arlock),               //  output,    width = 2,                   .arlock
		.m_dest_axi_rid     (axi_ad9680_dma_m_dest_axi_rid),                  //   input,    width = 1,                   .rid
		.m_dest_axi_bid     (axi_ad9680_dma_m_dest_axi_bid),                  //   input,    width = 1,                   .bid
		.m_dest_axi_rlast   (axi_ad9680_dma_m_dest_axi_rlast)                 //   input,    width = 1,                   .rlast
	);

	system_bd_sys_clk sys_clk (
		.in_clk      (sys_clk_clk),             //   input,  width = 1,       clk_in.clk
		.reset_n     (sys_rst_reset_n),         //   input,  width = 1, clk_in_reset.reset_n
		.clk_out     (sys_clk_clk_clk),         //  output,  width = 1,          clk.clk
		.reset_n_out (sys_clk_clk_reset_reset)  //  output,  width = 1,    clk_reset.reset_n
	);

	system_bd_sys_cpu sys_cpu (
		.clk                                 (sys_clk_clk_clk),                                       //   input,   width = 1,                                  clk.clk
		.reset_n                             (~rst_controller_004_reset_out_reset),                   //   input,   width = 1,                                reset.reset_n
		.reset_req                           (rst_controller_004_reset_out_reset_req),                //   input,   width = 1,                                     .reset_req
		.d_address                           (sys_cpu_data_master_address),                           //  output,  width = 29,                          data_master.address
		.d_byteenable                        (sys_cpu_data_master_byteenable),                        //  output,   width = 4,                                     .byteenable
		.d_read                              (sys_cpu_data_master_read),                              //  output,   width = 1,                                     .read
		.d_readdata                          (sys_cpu_data_master_readdata),                          //   input,  width = 32,                                     .readdata
		.d_waitrequest                       (sys_cpu_data_master_waitrequest),                       //   input,   width = 1,                                     .waitrequest
		.d_write                             (sys_cpu_data_master_write),                             //  output,   width = 1,                                     .write
		.d_writedata                         (sys_cpu_data_master_writedata),                         //  output,  width = 32,                                     .writedata
		.d_readdatavalid                     (sys_cpu_data_master_readdatavalid),                     //   input,   width = 1,                                     .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (sys_cpu_data_master_debugaccess),                       //  output,   width = 1,                                     .debugaccess
		.i_address                           (sys_cpu_instruction_master_address),                    //  output,  width = 29,                   instruction_master.address
		.i_read                              (sys_cpu_instruction_master_read),                       //  output,   width = 1,                                     .read
		.i_readdata                          (sys_cpu_instruction_master_readdata),                   //   input,  width = 32,                                     .readdata
		.i_waitrequest                       (sys_cpu_instruction_master_waitrequest),                //   input,   width = 1,                                     .waitrequest
		.i_readdatavalid                     (sys_cpu_instruction_master_readdatavalid),              //   input,   width = 1,                                     .readdatavalid
		.dtcm0_readdata                      (sys_cpu_tightly_coupled_data_master_0_readdata),        //   input,  width = 32,        tightly_coupled_data_master_0.readdata
		.dtcm0_address                       (sys_cpu_tightly_coupled_data_master_0_address),         //  output,  width = 29,                                     .address
		.dtcm0_read                          (sys_cpu_tightly_coupled_data_master_0_read),            //  output,   width = 1,                                     .read
		.dtcm0_write                         (sys_cpu_tightly_coupled_data_master_0_write),           //  output,   width = 1,                                     .write
		.dtcm0_writedata                     (sys_cpu_tightly_coupled_data_master_0_writedata),       //  output,  width = 32,                                     .writedata
		.dtcm0_byteenable                    (sys_cpu_tightly_coupled_data_master_0_byteenable),      //  output,   width = 4,                                     .byteenable
		.itcm0_readdata                      (sys_cpu_tightly_coupled_instruction_master_0_readdata), //   input,  width = 32, tightly_coupled_instruction_master_0.readdata
		.itcm0_address                       (sys_cpu_tightly_coupled_instruction_master_0_address),  //  output,  width = 29,                                     .address
		.itcm0_read                          (sys_cpu_tightly_coupled_instruction_master_0_read),     //  output,   width = 1,                                     .read
		.irq                                 (sys_cpu_irq_irq),                                       //   input,  width = 32,                                  irq.irq
		.debug_reset_request                 (sys_cpu_debug_reset_request_reset),                     //  output,   width = 1,                  debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_sys_cpu_debug_mem_slave_address),     //   input,   width = 9,                      debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_sys_cpu_debug_mem_slave_byteenable),  //   input,   width = 4,                                     .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_sys_cpu_debug_mem_slave_debugaccess), //   input,   width = 1,                                     .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_sys_cpu_debug_mem_slave_read),        //   input,   width = 1,                                     .read
		.debug_mem_slave_readdata            (mm_interconnect_0_sys_cpu_debug_mem_slave_readdata),    //  output,  width = 32,                                     .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_sys_cpu_debug_mem_slave_waitrequest), //  output,   width = 1,                                     .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_sys_cpu_debug_mem_slave_write),       //   input,   width = 1,                                     .write
		.debug_mem_slave_writedata           (mm_interconnect_0_sys_cpu_debug_mem_slave_writedata),   //   input,  width = 32,                                     .writedata
		.dummy_ci_port                       ()                                                       //  output,   width = 1,            custom_instruction_master.readra
	);

	system_bd_sys_ddr3_cntrl sys_ddr3_cntrl (
		.global_reset_n      (sys_clk_clk_reset_reset),                                   //   input,    width = 1,   global_reset_n.reset_n
		.pll_ref_clk         (sys_ddr3_cntrl_pll_ref_clk_clk),                            //   input,    width = 1,      pll_ref_clk.clk
		.oct_rzqin           (sys_ddr3_cntrl_oct_oct_rzqin),                              //   input,    width = 1,              oct.oct_rzqin
		.mem_ck              (sys_ddr3_cntrl_mem_mem_ck),                                 //  output,    width = 1,              mem.mem_ck
		.mem_ck_n            (sys_ddr3_cntrl_mem_mem_ck_n),                               //  output,    width = 1,                 .mem_ck_n
		.mem_a               (sys_ddr3_cntrl_mem_mem_a),                                  //  output,   width = 12,                 .mem_a
		.mem_ba              (sys_ddr3_cntrl_mem_mem_ba),                                 //  output,    width = 3,                 .mem_ba
		.mem_cke             (sys_ddr3_cntrl_mem_mem_cke),                                //  output,    width = 1,                 .mem_cke
		.mem_cs_n            (sys_ddr3_cntrl_mem_mem_cs_n),                               //  output,    width = 1,                 .mem_cs_n
		.mem_odt             (sys_ddr3_cntrl_mem_mem_odt),                                //  output,    width = 1,                 .mem_odt
		.mem_reset_n         (sys_ddr3_cntrl_mem_mem_reset_n),                            //  output,    width = 1,                 .mem_reset_n
		.mem_we_n            (sys_ddr3_cntrl_mem_mem_we_n),                               //  output,    width = 1,                 .mem_we_n
		.mem_ras_n           (sys_ddr3_cntrl_mem_mem_ras_n),                              //  output,    width = 1,                 .mem_ras_n
		.mem_cas_n           (sys_ddr3_cntrl_mem_mem_cas_n),                              //  output,    width = 1,                 .mem_cas_n
		.mem_dqs             (sys_ddr3_cntrl_mem_mem_dqs),                                //   inout,    width = 8,                 .mem_dqs
		.mem_dqs_n           (sys_ddr3_cntrl_mem_mem_dqs_n),                              //   inout,    width = 8,                 .mem_dqs_n
		.mem_dq              (sys_ddr3_cntrl_mem_mem_dq),                                 //   inout,   width = 64,                 .mem_dq
		.mem_dm              (sys_ddr3_cntrl_mem_mem_dm),                                 //  output,    width = 8,                 .mem_dm
		.local_cal_success   (),                                                          //  output,    width = 1,           status.local_cal_success
		.local_cal_fail      (),                                                          //  output,    width = 1,                 .local_cal_fail
		.emif_usr_reset_n    (sys_ddr3_cntrl_emif_usr_reset_n_reset),                     //  output,    width = 1, emif_usr_reset_n.reset_n
		.emif_usr_clk        (sys_ddr3_cntrl_emif_usr_clk_clk),                           //  output,    width = 1,     emif_usr_clk.clk
		.amm_ready_0         (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_waitrequest),   //  output,    width = 1,       ctrl_amm_0.waitrequest_n
		.amm_read_0          (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_read),          //   input,    width = 1,                 .read
		.amm_write_0         (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_write),         //   input,    width = 1,                 .write
		.amm_address_0       (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_address),       //   input,   width = 22,                 .address
		.amm_readdata_0      (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_readdata),      //  output,  width = 512,                 .readdata
		.amm_writedata_0     (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_writedata),     //   input,  width = 512,                 .writedata
		.amm_burstcount_0    (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_burstcount),    //   input,    width = 7,                 .burstcount
		.amm_byteenable_0    (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_byteenable),    //   input,   width = 64,                 .byteenable
		.amm_readdatavalid_0 (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_readdatavalid)  //  output,    width = 1,                 .readdatavalid
	);

	system_bd_sys_dma_clk sys_dma_clk (
		.in_clk      (sys_ddr3_cntrl_emif_usr_clk_clk),       //   input,  width = 1,       clk_in.clk
		.reset_n     (sys_ddr3_cntrl_emif_usr_reset_n_reset), //   input,  width = 1, clk_in_reset.reset_n
		.clk_out     (sys_dma_clk_clk_clk),                   //  output,  width = 1,          clk.clk
		.reset_n_out (sys_dma_clk_clk_reset_reset)            //  output,  width = 1,    clk_reset.reset_n
	);

	system_bd_sys_ethernet sys_ethernet (
		.ff_tx_clk      (sys_clk_clk_clk),                                         //   input,   width = 1,     transmit_clock_connection.clk
		.ff_rx_clk      (sys_clk_clk_clk),                                         //   input,   width = 1,      receive_clock_connection.clk
		.ff_rx_data     (sys_ethernet_receive_data),                               //  output,  width = 32,                       receive.data
		.ff_rx_eop      (sys_ethernet_receive_endofpacket),                        //  output,   width = 1,                              .endofpacket
		.rx_err         (sys_ethernet_receive_error),                              //  output,   width = 6,                              .error
		.ff_rx_mod      (sys_ethernet_receive_empty),                              //  output,   width = 2,                              .empty
		.ff_rx_rdy      (sys_ethernet_receive_ready),                              //   input,   width = 1,                              .ready
		.ff_rx_sop      (sys_ethernet_receive_startofpacket),                      //  output,   width = 1,                              .startofpacket
		.ff_rx_dval     (sys_ethernet_receive_valid),                              //  output,   width = 1,                              .valid
		.ff_tx_data     (avalon_st_adapter_001_out_0_data),                        //   input,  width = 32,                      transmit.data
		.ff_tx_eop      (avalon_st_adapter_001_out_0_endofpacket),                 //   input,   width = 1,                              .endofpacket
		.ff_tx_err      (avalon_st_adapter_001_out_0_error),                       //   input,   width = 1,                              .error
		.ff_tx_mod      (avalon_st_adapter_001_out_0_empty),                       //   input,   width = 2,                              .empty
		.ff_tx_rdy      (avalon_st_adapter_001_out_0_ready),                       //  output,   width = 1,                              .ready
		.ff_tx_sop      (avalon_st_adapter_001_out_0_startofpacket),               //   input,   width = 1,                              .startofpacket
		.ff_tx_wren     (avalon_st_adapter_001_out_0_valid),                       //   input,   width = 1,                              .valid
		.magic_wakeup   (),                                                        //  output,   width = 1,           mac_misc_connection.magic_wakeup
		.magic_sleep_n  (),                                                        //   input,   width = 1,                              .magic_sleep_n
		.ff_tx_crc_fwd  (),                                                        //   input,   width = 1,                              .ff_tx_crc_fwd
		.ff_tx_septy    (),                                                        //  output,   width = 1,                              .ff_tx_septy
		.tx_ff_uflow    (),                                                        //  output,   width = 1,                              .tx_ff_uflow
		.ff_tx_a_full   (),                                                        //  output,   width = 1,                              .ff_tx_a_full
		.ff_tx_a_empty  (),                                                        //  output,   width = 1,                              .ff_tx_a_empty
		.rx_err_stat    (),                                                        //  output,  width = 18,                              .rx_err_stat
		.rx_frm_type    (),                                                        //  output,   width = 4,                              .rx_frm_type
		.ff_rx_dsav     (),                                                        //  output,   width = 1,                              .ff_rx_dsav
		.ff_rx_a_full   (),                                                        //  output,   width = 1,                              .ff_rx_a_full
		.ff_rx_a_empty  (),                                                        //  output,   width = 1,                              .ff_rx_a_empty
		.mdc            (sys_ethernet_mdio_mdc),                                   //  output,   width = 1,           mac_mdio_connection.mdc
		.mdio_in        (sys_ethernet_mdio_mdio_in),                               //   input,   width = 1,                              .mdio_in
		.mdio_out       (sys_ethernet_mdio_mdio_out),                              //  output,   width = 1,                              .mdio_out
		.mdio_oen       (sys_ethernet_mdio_mdio_oen),                              //  output,   width = 1,                              .mdio_oen
		.clk            (sys_clk_clk_clk),                                         //   input,   width = 1, control_port_clock_connection.clk
		.reset          (rst_controller_reset_out_reset),                          //   input,   width = 1,              reset_connection.reset
		.reg_data_out   (mm_interconnect_0_sys_ethernet_control_port_readdata),    //  output,  width = 32,                  control_port.readdata
		.reg_rd         (mm_interconnect_0_sys_ethernet_control_port_read),        //   input,   width = 1,                              .read
		.reg_data_in    (mm_interconnect_0_sys_ethernet_control_port_writedata),   //   input,  width = 32,                              .writedata
		.reg_wr         (mm_interconnect_0_sys_ethernet_control_port_write),       //   input,   width = 1,                              .write
		.reg_busy       (mm_interconnect_0_sys_ethernet_control_port_waitrequest), //  output,   width = 1,                              .waitrequest
		.reg_addr       (mm_interconnect_0_sys_ethernet_control_port_address),     //   input,   width = 8,                              .address
		.ref_clk        (sys_ethernet_ref_clk_clk),                                //   input,   width = 1,  pcs_ref_clk_clock_connection.clk
		.led_crs        (),                                                        //  output,   width = 1,         status_led_connection.crs
		.led_link       (),                                                        //  output,   width = 1,                              .link
		.led_panel_link (),                                                        //  output,   width = 1,                              .panel_link
		.led_col        (),                                                        //  output,   width = 1,                              .col
		.led_an         (),                                                        //  output,   width = 1,                              .an
		.led_char_err   (),                                                        //  output,   width = 1,                              .char_err
		.led_disp_err   (),                                                        //  output,   width = 1,                              .disp_err
		.rx_recovclkout (),                                                        //  output,   width = 1,     serdes_control_connection.export
		.rxp            (sys_ethernet_sgmii_rxp_0),                                //   input,   width = 1,             serial_connection.rxp_0
		.txp            (sys_ethernet_sgmii_txp_0)                                 //  output,   width = 1,                              .txp_0
	);

	system_bd_sys_ethernet_dma_rx sys_ethernet_dma_rx (
		.clock_clk                    (sys_clk_clk_clk),                                                    //   input,    width = 1,            clock.clk
		.reset_n_reset_n              (~rst_controller_005_reset_out_reset),                                //   input,    width = 1,          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_sys_ethernet_dma_rx_csr_writedata),                //   input,   width = 32,              csr.writedata
		.csr_write                    (mm_interconnect_0_sys_ethernet_dma_rx_csr_write),                    //   input,    width = 1,                 .write
		.csr_byteenable               (mm_interconnect_0_sys_ethernet_dma_rx_csr_byteenable),               //   input,    width = 4,                 .byteenable
		.csr_readdata                 (mm_interconnect_0_sys_ethernet_dma_rx_csr_readdata),                 //  output,   width = 32,                 .readdata
		.csr_read                     (mm_interconnect_0_sys_ethernet_dma_rx_csr_read),                     //   input,    width = 1,                 .read
		.csr_address                  (mm_interconnect_0_sys_ethernet_dma_rx_csr_address),                  //   input,    width = 3,                 .address
		.descriptor_slave_write       (mm_interconnect_0_sys_ethernet_dma_rx_descriptor_slave_write),       //   input,    width = 1, descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_sys_ethernet_dma_rx_descriptor_slave_waitrequest), //  output,    width = 1,                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_sys_ethernet_dma_rx_descriptor_slave_writedata),   //   input,  width = 256,                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_sys_ethernet_dma_rx_descriptor_slave_byteenable),  //   input,   width = 32,                 .byteenable
		.response_waitrequest         (mm_interconnect_0_sys_ethernet_dma_rx_response_waitrequest),         //  output,    width = 1,         response.waitrequest
		.response_byteenable          (mm_interconnect_0_sys_ethernet_dma_rx_response_byteenable),          //   input,    width = 4,                 .byteenable
		.response_address             (mm_interconnect_0_sys_ethernet_dma_rx_response_address),             //   input,    width = 1,                 .address
		.response_readdata            (mm_interconnect_0_sys_ethernet_dma_rx_response_readdata),            //  output,   width = 32,                 .readdata
		.response_read                (mm_interconnect_0_sys_ethernet_dma_rx_response_read),                //   input,    width = 1,                 .read
		.csr_irq_irq                  (irq_mapper_receiver0_irq),                                           //  output,    width = 1,          csr_irq.irq
		.mm_write_address             (sys_ethernet_dma_rx_mm_write_address),                               //  output,   width = 32,         mm_write.address
		.mm_write_write               (sys_ethernet_dma_rx_mm_write_write),                                 //  output,    width = 1,                 .write
		.mm_write_byteenable          (sys_ethernet_dma_rx_mm_write_byteenable),                            //  output,    width = 8,                 .byteenable
		.mm_write_writedata           (sys_ethernet_dma_rx_mm_write_writedata),                             //  output,   width = 64,                 .writedata
		.mm_write_waitrequest         (sys_ethernet_dma_rx_mm_write_waitrequest),                           //   input,    width = 1,                 .waitrequest
		.mm_write_burstcount          (sys_ethernet_dma_rx_mm_write_burstcount),                            //  output,    width = 7,                 .burstcount
		.st_sink_data                 (avalon_st_adapter_out_0_data),                                       //   input,   width = 64,          st_sink.data
		.st_sink_valid                (avalon_st_adapter_out_0_valid),                                      //   input,    width = 1,                 .valid
		.st_sink_ready                (avalon_st_adapter_out_0_ready),                                      //  output,    width = 1,                 .ready
		.st_sink_startofpacket        (avalon_st_adapter_out_0_startofpacket),                              //   input,    width = 1,                 .startofpacket
		.st_sink_endofpacket          (avalon_st_adapter_out_0_endofpacket),                                //   input,    width = 1,                 .endofpacket
		.st_sink_empty                (avalon_st_adapter_out_0_empty),                                      //   input,    width = 3,                 .empty
		.st_sink_error                (avalon_st_adapter_out_0_error)                                       //   input,    width = 6,                 .error
	);

	system_bd_sys_ethernet_dma_tx sys_ethernet_dma_tx (
		.clock_clk                    (sys_clk_clk_clk),                                                    //   input,    width = 1,            clock.clk
		.reset_n_reset_n              (~rst_controller_005_reset_out_reset),                                //   input,    width = 1,          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_sys_ethernet_dma_tx_csr_writedata),                //   input,   width = 32,              csr.writedata
		.csr_write                    (mm_interconnect_0_sys_ethernet_dma_tx_csr_write),                    //   input,    width = 1,                 .write
		.csr_byteenable               (mm_interconnect_0_sys_ethernet_dma_tx_csr_byteenable),               //   input,    width = 4,                 .byteenable
		.csr_readdata                 (mm_interconnect_0_sys_ethernet_dma_tx_csr_readdata),                 //  output,   width = 32,                 .readdata
		.csr_read                     (mm_interconnect_0_sys_ethernet_dma_tx_csr_read),                     //   input,    width = 1,                 .read
		.csr_address                  (mm_interconnect_0_sys_ethernet_dma_tx_csr_address),                  //   input,    width = 3,                 .address
		.descriptor_slave_write       (mm_interconnect_0_sys_ethernet_dma_tx_descriptor_slave_write),       //   input,    width = 1, descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_sys_ethernet_dma_tx_descriptor_slave_waitrequest), //  output,    width = 1,                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_sys_ethernet_dma_tx_descriptor_slave_writedata),   //   input,  width = 256,                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_sys_ethernet_dma_tx_descriptor_slave_byteenable),  //   input,   width = 32,                 .byteenable
		.csr_irq_irq                  (irq_mapper_receiver1_irq),                                           //  output,    width = 1,          csr_irq.irq
		.mm_read_address              (sys_ethernet_dma_tx_mm_read_address),                                //  output,   width = 32,          mm_read.address
		.mm_read_read                 (sys_ethernet_dma_tx_mm_read_read),                                   //  output,    width = 1,                 .read
		.mm_read_byteenable           (sys_ethernet_dma_tx_mm_read_byteenable),                             //  output,    width = 8,                 .byteenable
		.mm_read_readdata             (sys_ethernet_dma_tx_mm_read_readdata),                               //   input,   width = 64,                 .readdata
		.mm_read_waitrequest          (sys_ethernet_dma_tx_mm_read_waitrequest),                            //   input,    width = 1,                 .waitrequest
		.mm_read_readdatavalid        (sys_ethernet_dma_tx_mm_read_readdatavalid),                          //   input,    width = 1,                 .readdatavalid
		.mm_read_burstcount           (sys_ethernet_dma_tx_mm_read_burstcount),                             //  output,    width = 7,                 .burstcount
		.st_source_data               (sys_ethernet_dma_tx_st_source_data),                                 //  output,   width = 64,        st_source.data
		.st_source_valid              (sys_ethernet_dma_tx_st_source_valid),                                //  output,    width = 1,                 .valid
		.st_source_ready              (sys_ethernet_dma_tx_st_source_ready),                                //   input,    width = 1,                 .ready
		.st_source_startofpacket      (sys_ethernet_dma_tx_st_source_startofpacket),                        //  output,    width = 1,                 .startofpacket
		.st_source_endofpacket        (sys_ethernet_dma_tx_st_source_endofpacket),                          //  output,    width = 1,                 .endofpacket
		.st_source_empty              (sys_ethernet_dma_tx_st_source_empty),                                //  output,    width = 3,                 .empty
		.st_source_error              (sys_ethernet_dma_tx_st_source_error)                                 //  output,    width = 1,                 .error
	);

	system_bd_sys_ethernet_reset sys_ethernet_reset (
		.clk       (sys_clk_clk_clk),                //   input,  width = 1,       clk.clk
		.in_reset  (rst_controller_reset_out_reset), //   input,  width = 1,  in_reset.reset
		.out_reset (sys_ethernet_reset_reset)        //  output,  width = 1, out_reset.reset
	);

	system_bd_sys_flash sys_flash (
		.clk_clk              (sys_clk_clk_clk),                               //   input,   width = 1,   clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                //   input,   width = 1, reset.reset
		.uas_address          (mm_interconnect_0_sys_flash_uas_address),       //   input,  width = 24,   uas.address
		.uas_burstcount       (mm_interconnect_0_sys_flash_uas_burstcount),    //   input,   width = 3,      .burstcount
		.uas_read             (mm_interconnect_0_sys_flash_uas_read),          //   input,   width = 1,      .read
		.uas_write            (mm_interconnect_0_sys_flash_uas_write),         //   input,   width = 1,      .write
		.uas_waitrequest      (mm_interconnect_0_sys_flash_uas_waitrequest),   //  output,   width = 1,      .waitrequest
		.uas_readdatavalid    (mm_interconnect_0_sys_flash_uas_readdatavalid), //  output,   width = 1,      .readdatavalid
		.uas_byteenable       (mm_interconnect_0_sys_flash_uas_byteenable),    //   input,   width = 4,      .byteenable
		.uas_readdata         (mm_interconnect_0_sys_flash_uas_readdata),      //  output,  width = 32,      .readdata
		.uas_writedata        (mm_interconnect_0_sys_flash_uas_writedata),     //   input,  width = 32,      .writedata
		.uas_lock             (mm_interconnect_0_sys_flash_uas_lock),          //   input,   width = 1,      .lock
		.uas_debugaccess      (mm_interconnect_0_sys_flash_uas_debugaccess),   //   input,   width = 1,      .debugaccess
		.tcm_write_n_out      (sys_flash_tcm_write_n_out_signal),              //  output,   width = 1,   tcm.write_n_out
		.tcm_read_n_out       (sys_flash_tcm_read_n_out_signal),               //  output,   width = 1,      .read_n_out
		.tcm_chipselect_n_out (sys_flash_tcm_chipselect_n_out_signal),         //  output,   width = 1,      .chipselect_n_out
		.tcm_request          (sys_flash_tcm_request),                         //  output,   width = 1,      .request
		.tcm_grant            (sys_flash_tcm_grant),                           //   input,   width = 1,      .grant
		.tcm_address_out      (sys_flash_tcm_address_out_signal),              //  output,  width = 24,      .address_out
		.tcm_data_out         (sys_flash_tcm_data_out_signal),                 //  output,  width = 32,      .data_out
		.tcm_data_outen       (sys_flash_tcm_data_outen),                      //  output,   width = 1,      .data_outen
		.tcm_data_in          (sys_flash_tcm_data_in)                          //   input,  width = 32,      .data_in
	);

	system_bd_sys_flash_bridge sys_flash_bridge (
		.clk                      (sys_clk_clk_clk),                       //   input,   width = 1,   clk.clk
		.reset                    (rst_controller_reset_out_reset),        //   input,   width = 1, reset.reset
		.request                  (sys_flash_tcm_request),                 //   input,   width = 1,   tcs.request
		.grant                    (sys_flash_tcm_grant),                   //  output,   width = 1,      .grant
		.tcs_tcm_address_out      (sys_flash_tcm_address_out_signal),      //   input,  width = 24,      .address_out
		.tcs_tcm_read_n_out       (sys_flash_tcm_read_n_out_signal),       //   input,   width = 1,      .read_n_out
		.tcs_tcm_write_n_out      (sys_flash_tcm_write_n_out_signal),      //   input,   width = 1,      .write_n_out
		.tcs_tcm_data_out         (sys_flash_tcm_data_out_signal),         //   input,  width = 32,      .data_out
		.tcs_tcm_data_outen       (sys_flash_tcm_data_outen),              //   input,   width = 1,      .data_outen
		.tcs_tcm_data_in          (sys_flash_tcm_data_in),                 //  output,  width = 32,      .data_in
		.tcs_tcm_chipselect_n_out (sys_flash_tcm_chipselect_n_out_signal), //   input,   width = 1,      .chipselect_n_out
		.tcm_address_out          (sys_flash_tcm_address_out),             //  output,  width = 24,   out.tcm_address_out
		.tcm_read_n_out           (sys_flash_tcm_read_n_out),              //  output,   width = 1,      .tcm_read_n_out
		.tcm_write_n_out          (sys_flash_tcm_write_n_out),             //  output,   width = 1,      .tcm_write_n_out
		.tcm_data_out             (sys_flash_tcm_data_out),                //   inout,  width = 32,      .tcm_data_out
		.tcm_chipselect_n_out     (sys_flash_tcm_chipselect_n_out)         //  output,   width = 1,      .tcm_chipselect_n_out
	);

	system_bd_sys_gpio_bd sys_gpio_bd (
		.clk        (sys_clk_clk_clk),                             //   input,   width = 1,                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //   input,   width = 1,               reset.reset_n
		.address    (mm_interconnect_0_sys_gpio_bd_s1_address),    //   input,   width = 2,                  s1.address
		.write_n    (~mm_interconnect_0_sys_gpio_bd_s1_write),     //   input,   width = 1,                    .write_n
		.writedata  (mm_interconnect_0_sys_gpio_bd_s1_writedata),  //   input,  width = 32,                    .writedata
		.chipselect (mm_interconnect_0_sys_gpio_bd_s1_chipselect), //   input,   width = 1,                    .chipselect
		.readdata   (mm_interconnect_0_sys_gpio_bd_s1_readdata),   //  output,  width = 32,                    .readdata
		.in_port    (sys_gpio_bd_in_port),                         //   input,  width = 32, external_connection.in_port
		.out_port   (sys_gpio_bd_out_port),                        //  output,  width = 32,                    .out_port
		.irq        (irq_mapper_receiver8_irq)                     //  output,   width = 1,                 irq.irq
	);

	system_bd_sys_gpio_in sys_gpio_in (
		.clk        (sys_clk_clk_clk),                             //   input,   width = 1,                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //   input,   width = 1,               reset.reset_n
		.address    (mm_interconnect_0_sys_gpio_in_s1_address),    //   input,   width = 2,                  s1.address
		.write_n    (~mm_interconnect_0_sys_gpio_in_s1_write),     //   input,   width = 1,                    .write_n
		.writedata  (mm_interconnect_0_sys_gpio_in_s1_writedata),  //   input,  width = 32,                    .writedata
		.chipselect (mm_interconnect_0_sys_gpio_in_s1_chipselect), //   input,   width = 1,                    .chipselect
		.readdata   (mm_interconnect_0_sys_gpio_in_s1_readdata),   //  output,  width = 32,                    .readdata
		.in_port    (sys_gpio_in_export),                          //   input,  width = 32, external_connection.export
		.irq        (irq_mapper_receiver7_irq)                     //  output,   width = 1,                 irq.irq
	);

	system_bd_sys_gpio_out sys_gpio_out (
		.clk        (sys_clk_clk_clk),                              //   input,   width = 1,                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //   input,   width = 1,               reset.reset_n
		.address    (mm_interconnect_0_sys_gpio_out_s1_address),    //   input,   width = 2,                  s1.address
		.write_n    (~mm_interconnect_0_sys_gpio_out_s1_write),     //   input,   width = 1,                    .write_n
		.writedata  (mm_interconnect_0_sys_gpio_out_s1_writedata),  //   input,  width = 32,                    .writedata
		.chipselect (mm_interconnect_0_sys_gpio_out_s1_chipselect), //   input,   width = 1,                    .chipselect
		.readdata   (mm_interconnect_0_sys_gpio_out_s1_readdata),   //  output,  width = 32,                    .readdata
		.out_port   (sys_gpio_out_export)                           //  output,  width = 32, external_connection.export
	);

	system_bd_sys_id sys_id (
		.clock    (sys_clk_clk_clk),                                 //   input,   width = 1,           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //   input,   width = 1,         reset.reset_n
		.readdata (mm_interconnect_0_sys_id_control_slave_readdata), //  output,  width = 32, control_slave.readdata
		.address  (mm_interconnect_0_sys_id_control_slave_address)   //   input,   width = 1,              .address
	);

	system_bd_sys_int_mem sys_int_mem (
		.clk        (sys_clk_clk_clk),                             //   input,   width = 1,   clk1.clk
		.address    (mm_interconnect_0_sys_int_mem_s1_address),    //   input,  width = 16,     s1.address
		.clken      (mm_interconnect_0_sys_int_mem_s1_clken),      //   input,   width = 1,       .clken
		.chipselect (mm_interconnect_0_sys_int_mem_s1_chipselect), //   input,   width = 1,       .chipselect
		.write      (mm_interconnect_0_sys_int_mem_s1_write),      //   input,   width = 1,       .write
		.readdata   (mm_interconnect_0_sys_int_mem_s1_readdata),   //  output,  width = 32,       .readdata
		.writedata  (mm_interconnect_0_sys_int_mem_s1_writedata),  //   input,  width = 32,       .writedata
		.byteenable (mm_interconnect_0_sys_int_mem_s1_byteenable), //   input,   width = 4,       .byteenable
		.reset      (rst_controller_reset_out_reset),              //   input,   width = 1, reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)           //   input,   width = 1,       .reset_req
	);

	system_bd_sys_spi sys_spi (
		.clk           (sys_clk_clk_clk),                                       //   input,   width = 1,              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //   input,   width = 1,            reset.reset_n
		.data_from_cpu (mm_interconnect_0_sys_spi_spi_control_port_writedata),  //   input,  width = 16, spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_sys_spi_spi_control_port_readdata),   //  output,  width = 16,                 .readdata
		.mem_addr      (mm_interconnect_0_sys_spi_spi_control_port_address),    //   input,   width = 3,                 .address
		.read_n        (~mm_interconnect_0_sys_spi_spi_control_port_read),      //   input,   width = 1,                 .read_n
		.spi_select    (mm_interconnect_0_sys_spi_spi_control_port_chipselect), //   input,   width = 1,                 .chipselect
		.write_n       (~mm_interconnect_0_sys_spi_spi_control_port_write),     //   input,   width = 1,                 .write_n
		.irq           (irq_mapper_receiver9_irq),                              //  output,   width = 1,              irq.irq
		.MISO          (sys_spi_MISO),                                          //   input,   width = 1,         external.MISO
		.MOSI          (sys_spi_MOSI),                                          //  output,   width = 1,                 .MOSI
		.SCLK          (sys_spi_SCLK),                                          //  output,   width = 1,                 .SCLK
		.SS_n          (sys_spi_SS_n)                                           //  output,   width = 8,                 .SS_n
	);

	system_bd_sys_timer_1 sys_timer_1 (
		.clk        (sys_clk_clk_clk),                             //   input,   width = 1,   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //   input,   width = 1, reset.reset_n
		.address    (mm_interconnect_0_sys_timer_1_s1_address),    //   input,   width = 3,    s1.address
		.writedata  (mm_interconnect_0_sys_timer_1_s1_writedata),  //   input,  width = 16,      .writedata
		.readdata   (mm_interconnect_0_sys_timer_1_s1_readdata),   //  output,  width = 16,      .readdata
		.chipselect (mm_interconnect_0_sys_timer_1_s1_chipselect), //   input,   width = 1,      .chipselect
		.write_n    (~mm_interconnect_0_sys_timer_1_s1_write),     //   input,   width = 1,      .write_n
		.irq        (irq_mapper_receiver6_irq)                     //  output,   width = 1,   irq.irq
	);

	system_bd_sys_timer_2 sys_timer_2 (
		.clk        (sys_clk_clk_clk),                             //   input,   width = 1,   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //   input,   width = 1, reset.reset_n
		.address    (mm_interconnect_0_sys_timer_2_s1_address),    //   input,   width = 3,    s1.address
		.writedata  (mm_interconnect_0_sys_timer_2_s1_writedata),  //   input,  width = 16,      .writedata
		.readdata   (mm_interconnect_0_sys_timer_2_s1_readdata),   //  output,  width = 16,      .readdata
		.chipselect (mm_interconnect_0_sys_timer_2_s1_chipselect), //   input,   width = 1,      .chipselect
		.write_n    (~mm_interconnect_0_sys_timer_2_s1_write),     //   input,   width = 1,      .write_n
		.irq        (irq_mapper_receiver5_irq)                     //  output,   width = 1,   irq.irq
	);

	system_bd_sys_tlb_mem sys_tlb_mem (
		.clk         (sys_clk_clk_clk),                             //   input,   width = 1,   clk1.clk
		.address     (mm_interconnect_1_sys_tlb_mem_s1_address),    //   input,  width = 16,     s1.address
		.clken       (mm_interconnect_1_sys_tlb_mem_s1_clken),      //   input,   width = 1,       .clken
		.chipselect  (mm_interconnect_1_sys_tlb_mem_s1_chipselect), //   input,   width = 1,       .chipselect
		.write       (mm_interconnect_1_sys_tlb_mem_s1_write),      //   input,   width = 1,       .write
		.readdata    (mm_interconnect_1_sys_tlb_mem_s1_readdata),   //  output,  width = 32,       .readdata
		.writedata   (mm_interconnect_1_sys_tlb_mem_s1_writedata),  //   input,  width = 32,       .writedata
		.byteenable  (mm_interconnect_1_sys_tlb_mem_s1_byteenable), //   input,   width = 4,       .byteenable
		.reset       (rst_controller_reset_out_reset),              //   input,   width = 1, reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //   input,   width = 1,       .reset_req
		.address2    (mm_interconnect_2_sys_tlb_mem_s2_address),    //   input,  width = 16,     s2.address
		.chipselect2 (mm_interconnect_2_sys_tlb_mem_s2_chipselect), //   input,   width = 1,       .chipselect
		.clken2      (mm_interconnect_2_sys_tlb_mem_s2_clken),      //   input,   width = 1,       .clken
		.write2      (mm_interconnect_2_sys_tlb_mem_s2_write),      //   input,   width = 1,       .write
		.readdata2   (mm_interconnect_2_sys_tlb_mem_s2_readdata),   //  output,  width = 32,       .readdata
		.writedata2  (mm_interconnect_2_sys_tlb_mem_s2_writedata),  //   input,  width = 32,       .writedata
		.byteenable2 (mm_interconnect_2_sys_tlb_mem_s2_byteenable), //   input,   width = 4,       .byteenable
		.clk2        (sys_clk_clk_clk),                             //   input,   width = 1,   clk2.clk
		.reset2      (rst_controller_reset_out_reset),              //   input,   width = 1, reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req)           //   input,   width = 1,       .reset_req
	);

	system_bd_sys_uart sys_uart (
		.clk            (sys_clk_clk_clk),                                          //   input,   width = 1,               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                          //   input,   width = 1,             reset.reset_n
		.av_chipselect  (mm_interconnect_0_sys_uart_avalon_jtag_slave_chipselect),  //   input,   width = 1, avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_sys_uart_avalon_jtag_slave_address),     //   input,   width = 1,                  .address
		.av_read_n      (~mm_interconnect_0_sys_uart_avalon_jtag_slave_read),       //   input,   width = 1,                  .read_n
		.av_readdata    (mm_interconnect_0_sys_uart_avalon_jtag_slave_readdata),    //  output,  width = 32,                  .readdata
		.av_write_n     (~mm_interconnect_0_sys_uart_avalon_jtag_slave_write),      //   input,   width = 1,                  .write_n
		.av_writedata   (mm_interconnect_0_sys_uart_avalon_jtag_slave_writedata),   //   input,  width = 32,                  .writedata
		.av_waitrequest (mm_interconnect_0_sys_uart_avalon_jtag_slave_waitrequest), //  output,   width = 1,                  .waitrequest
		.av_irq         (irq_mapper_receiver4_irq)                                  //  output,   width = 1,               irq.irq
	);

	system_bd_util_ad9144_upack util_ad9144_upack (
		.dac_clk         (ad9144_jesd204_link_clk_clk),          //   input,    width = 1,   if_dac_clk.clk
		.dac_valid       (util_ad9144_upack_if_dac_valid_valid), //  output,    width = 1, if_dac_valid.valid
		.dac_sync        (),                                     //  output,    width = 1,  if_dac_sync.sync
		.dac_data        (avl_ad9144_fifo_if_dac_data_data),     //   input,  width = 128,  if_dac_data.data
		.dac_enable_0    (),                                     //   input,    width = 1,     dac_ch_0.enable
		.dac_valid_0     (),                                     //   input,    width = 1,             .valid
		.dac_valid_out_0 (),                                     //  output,    width = 1,             .data_valid
		.dac_data_0      (),                                     //  output,   width = 64,             .data
		.dac_enable_1    (),                                     //   input,    width = 1,     dac_ch_1.enable
		.dac_valid_1     (),                                     //   input,    width = 1,             .valid
		.dac_valid_out_1 (),                                     //  output,    width = 1,             .data_valid
		.dac_data_1      ()                                      //  output,   width = 64,             .data
	);

	system_bd_util_ad9680_cpack util_ad9680_cpack (
	);

	system_bd_altera_mm_interconnect_181_hkrcrsq mm_interconnect_0 (
		.sys_cpu_data_master_address                                            (sys_cpu_data_master_address),                                        //   input,   width = 29,                                              sys_cpu_data_master.address
		.sys_cpu_data_master_waitrequest                                        (sys_cpu_data_master_waitrequest),                                    //  output,    width = 1,                                                                 .waitrequest
		.sys_cpu_data_master_byteenable                                         (sys_cpu_data_master_byteenable),                                     //   input,    width = 4,                                                                 .byteenable
		.sys_cpu_data_master_read                                               (sys_cpu_data_master_read),                                           //   input,    width = 1,                                                                 .read
		.sys_cpu_data_master_readdata                                           (sys_cpu_data_master_readdata),                                       //  output,   width = 32,                                                                 .readdata
		.sys_cpu_data_master_readdatavalid                                      (sys_cpu_data_master_readdatavalid),                                  //  output,    width = 1,                                                                 .readdatavalid
		.sys_cpu_data_master_write                                              (sys_cpu_data_master_write),                                          //   input,    width = 1,                                                                 .write
		.sys_cpu_data_master_writedata                                          (sys_cpu_data_master_writedata),                                      //   input,   width = 32,                                                                 .writedata
		.sys_cpu_data_master_debugaccess                                        (sys_cpu_data_master_debugaccess),                                    //   input,    width = 1,                                                                 .debugaccess
		.sys_cpu_instruction_master_address                                     (sys_cpu_instruction_master_address),                                 //   input,   width = 29,                                       sys_cpu_instruction_master.address
		.sys_cpu_instruction_master_waitrequest                                 (sys_cpu_instruction_master_waitrequest),                             //  output,    width = 1,                                                                 .waitrequest
		.sys_cpu_instruction_master_read                                        (sys_cpu_instruction_master_read),                                    //   input,    width = 1,                                                                 .read
		.sys_cpu_instruction_master_readdata                                    (sys_cpu_instruction_master_readdata),                                //  output,   width = 32,                                                                 .readdata
		.sys_cpu_instruction_master_readdatavalid                               (sys_cpu_instruction_master_readdatavalid),                           //  output,    width = 1,                                                                 .readdatavalid
		.sys_ethernet_dma_tx_mm_read_address                                    (sys_ethernet_dma_tx_mm_read_address),                                //   input,   width = 32,                                      sys_ethernet_dma_tx_mm_read.address
		.sys_ethernet_dma_tx_mm_read_waitrequest                                (sys_ethernet_dma_tx_mm_read_waitrequest),                            //  output,    width = 1,                                                                 .waitrequest
		.sys_ethernet_dma_tx_mm_read_burstcount                                 (sys_ethernet_dma_tx_mm_read_burstcount),                             //   input,    width = 7,                                                                 .burstcount
		.sys_ethernet_dma_tx_mm_read_byteenable                                 (sys_ethernet_dma_tx_mm_read_byteenable),                             //   input,    width = 8,                                                                 .byteenable
		.sys_ethernet_dma_tx_mm_read_read                                       (sys_ethernet_dma_tx_mm_read_read),                                   //   input,    width = 1,                                                                 .read
		.sys_ethernet_dma_tx_mm_read_readdata                                   (sys_ethernet_dma_tx_mm_read_readdata),                               //  output,   width = 64,                                                                 .readdata
		.sys_ethernet_dma_tx_mm_read_readdatavalid                              (sys_ethernet_dma_tx_mm_read_readdatavalid),                          //  output,    width = 1,                                                                 .readdatavalid
		.sys_ethernet_dma_rx_mm_write_address                                   (sys_ethernet_dma_rx_mm_write_address),                               //   input,   width = 32,                                     sys_ethernet_dma_rx_mm_write.address
		.sys_ethernet_dma_rx_mm_write_waitrequest                               (sys_ethernet_dma_rx_mm_write_waitrequest),                           //  output,    width = 1,                                                                 .waitrequest
		.sys_ethernet_dma_rx_mm_write_burstcount                                (sys_ethernet_dma_rx_mm_write_burstcount),                            //   input,    width = 7,                                                                 .burstcount
		.sys_ethernet_dma_rx_mm_write_byteenable                                (sys_ethernet_dma_rx_mm_write_byteenable),                            //   input,    width = 8,                                                                 .byteenable
		.sys_ethernet_dma_rx_mm_write_write                                     (sys_ethernet_dma_rx_mm_write_write),                                 //   input,    width = 1,                                                                 .write
		.sys_ethernet_dma_rx_mm_write_writedata                                 (sys_ethernet_dma_rx_mm_write_writedata),                             //   input,   width = 64,                                                                 .writedata
		.sys_uart_avalon_jtag_slave_address                                     (mm_interconnect_0_sys_uart_avalon_jtag_slave_address),               //  output,    width = 1,                                       sys_uart_avalon_jtag_slave.address
		.sys_uart_avalon_jtag_slave_write                                       (mm_interconnect_0_sys_uart_avalon_jtag_slave_write),                 //  output,    width = 1,                                                                 .write
		.sys_uart_avalon_jtag_slave_read                                        (mm_interconnect_0_sys_uart_avalon_jtag_slave_read),                  //  output,    width = 1,                                                                 .read
		.sys_uart_avalon_jtag_slave_readdata                                    (mm_interconnect_0_sys_uart_avalon_jtag_slave_readdata),              //   input,   width = 32,                                                                 .readdata
		.sys_uart_avalon_jtag_slave_writedata                                   (mm_interconnect_0_sys_uart_avalon_jtag_slave_writedata),             //  output,   width = 32,                                                                 .writedata
		.sys_uart_avalon_jtag_slave_waitrequest                                 (mm_interconnect_0_sys_uart_avalon_jtag_slave_waitrequest),           //   input,    width = 1,                                                                 .waitrequest
		.sys_uart_avalon_jtag_slave_chipselect                                  (mm_interconnect_0_sys_uart_avalon_jtag_slave_chipselect),            //  output,    width = 1,                                                                 .chipselect
		.sys_ethernet_control_port_address                                      (mm_interconnect_0_sys_ethernet_control_port_address),                //  output,    width = 8,                                        sys_ethernet_control_port.address
		.sys_ethernet_control_port_write                                        (mm_interconnect_0_sys_ethernet_control_port_write),                  //  output,    width = 1,                                                                 .write
		.sys_ethernet_control_port_read                                         (mm_interconnect_0_sys_ethernet_control_port_read),                   //  output,    width = 1,                                                                 .read
		.sys_ethernet_control_port_readdata                                     (mm_interconnect_0_sys_ethernet_control_port_readdata),               //   input,   width = 32,                                                                 .readdata
		.sys_ethernet_control_port_writedata                                    (mm_interconnect_0_sys_ethernet_control_port_writedata),              //  output,   width = 32,                                                                 .writedata
		.sys_ethernet_control_port_waitrequest                                  (mm_interconnect_0_sys_ethernet_control_port_waitrequest),            //   input,    width = 1,                                                                 .waitrequest
		.sys_id_control_slave_address                                           (mm_interconnect_0_sys_id_control_slave_address),                     //  output,    width = 1,                                             sys_id_control_slave.address
		.sys_id_control_slave_readdata                                          (mm_interconnect_0_sys_id_control_slave_readdata),                    //   input,   width = 32,                                                                 .readdata
		.sys_ethernet_dma_rx_csr_address                                        (mm_interconnect_0_sys_ethernet_dma_rx_csr_address),                  //  output,    width = 3,                                          sys_ethernet_dma_rx_csr.address
		.sys_ethernet_dma_rx_csr_write                                          (mm_interconnect_0_sys_ethernet_dma_rx_csr_write),                    //  output,    width = 1,                                                                 .write
		.sys_ethernet_dma_rx_csr_read                                           (mm_interconnect_0_sys_ethernet_dma_rx_csr_read),                     //  output,    width = 1,                                                                 .read
		.sys_ethernet_dma_rx_csr_readdata                                       (mm_interconnect_0_sys_ethernet_dma_rx_csr_readdata),                 //   input,   width = 32,                                                                 .readdata
		.sys_ethernet_dma_rx_csr_writedata                                      (mm_interconnect_0_sys_ethernet_dma_rx_csr_writedata),                //  output,   width = 32,                                                                 .writedata
		.sys_ethernet_dma_rx_csr_byteenable                                     (mm_interconnect_0_sys_ethernet_dma_rx_csr_byteenable),               //  output,    width = 4,                                                                 .byteenable
		.sys_ethernet_dma_tx_csr_address                                        (mm_interconnect_0_sys_ethernet_dma_tx_csr_address),                  //  output,    width = 3,                                          sys_ethernet_dma_tx_csr.address
		.sys_ethernet_dma_tx_csr_write                                          (mm_interconnect_0_sys_ethernet_dma_tx_csr_write),                    //  output,    width = 1,                                                                 .write
		.sys_ethernet_dma_tx_csr_read                                           (mm_interconnect_0_sys_ethernet_dma_tx_csr_read),                     //  output,    width = 1,                                                                 .read
		.sys_ethernet_dma_tx_csr_readdata                                       (mm_interconnect_0_sys_ethernet_dma_tx_csr_readdata),                 //   input,   width = 32,                                                                 .readdata
		.sys_ethernet_dma_tx_csr_writedata                                      (mm_interconnect_0_sys_ethernet_dma_tx_csr_writedata),                //  output,   width = 32,                                                                 .writedata
		.sys_ethernet_dma_tx_csr_byteenable                                     (mm_interconnect_0_sys_ethernet_dma_tx_csr_byteenable),               //  output,    width = 4,                                                                 .byteenable
		.sys_ddr3_cntrl_ctrl_amm_0_address                                      (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_address),                //  output,   width = 22,                                        sys_ddr3_cntrl_ctrl_amm_0.address
		.sys_ddr3_cntrl_ctrl_amm_0_write                                        (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_write),                  //  output,    width = 1,                                                                 .write
		.sys_ddr3_cntrl_ctrl_amm_0_read                                         (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_read),                   //  output,    width = 1,                                                                 .read
		.sys_ddr3_cntrl_ctrl_amm_0_readdata                                     (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_readdata),               //   input,  width = 512,                                                                 .readdata
		.sys_ddr3_cntrl_ctrl_amm_0_writedata                                    (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_writedata),              //  output,  width = 512,                                                                 .writedata
		.sys_ddr3_cntrl_ctrl_amm_0_burstcount                                   (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_burstcount),             //  output,    width = 7,                                                                 .burstcount
		.sys_ddr3_cntrl_ctrl_amm_0_byteenable                                   (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_byteenable),             //  output,   width = 64,                                                                 .byteenable
		.sys_ddr3_cntrl_ctrl_amm_0_readdatavalid                                (mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_readdatavalid),          //   input,    width = 1,                                                                 .readdatavalid
		.sys_ddr3_cntrl_ctrl_amm_0_waitrequest                                  (~mm_interconnect_0_sys_ddr3_cntrl_ctrl_amm_0_waitrequest),           //   input,    width = 1,                                                                 .waitrequest
		.sys_cpu_debug_mem_slave_address                                        (mm_interconnect_0_sys_cpu_debug_mem_slave_address),                  //  output,    width = 9,                                          sys_cpu_debug_mem_slave.address
		.sys_cpu_debug_mem_slave_write                                          (mm_interconnect_0_sys_cpu_debug_mem_slave_write),                    //  output,    width = 1,                                                                 .write
		.sys_cpu_debug_mem_slave_read                                           (mm_interconnect_0_sys_cpu_debug_mem_slave_read),                     //  output,    width = 1,                                                                 .read
		.sys_cpu_debug_mem_slave_readdata                                       (mm_interconnect_0_sys_cpu_debug_mem_slave_readdata),                 //   input,   width = 32,                                                                 .readdata
		.sys_cpu_debug_mem_slave_writedata                                      (mm_interconnect_0_sys_cpu_debug_mem_slave_writedata),                //  output,   width = 32,                                                                 .writedata
		.sys_cpu_debug_mem_slave_byteenable                                     (mm_interconnect_0_sys_cpu_debug_mem_slave_byteenable),               //  output,    width = 4,                                                                 .byteenable
		.sys_cpu_debug_mem_slave_waitrequest                                    (mm_interconnect_0_sys_cpu_debug_mem_slave_waitrequest),              //   input,    width = 1,                                                                 .waitrequest
		.sys_cpu_debug_mem_slave_debugaccess                                    (mm_interconnect_0_sys_cpu_debug_mem_slave_debugaccess),              //  output,    width = 1,                                                                 .debugaccess
		.sys_ethernet_dma_rx_descriptor_slave_write                             (mm_interconnect_0_sys_ethernet_dma_rx_descriptor_slave_write),       //  output,    width = 1,                             sys_ethernet_dma_rx_descriptor_slave.write
		.sys_ethernet_dma_rx_descriptor_slave_writedata                         (mm_interconnect_0_sys_ethernet_dma_rx_descriptor_slave_writedata),   //  output,  width = 256,                                                                 .writedata
		.sys_ethernet_dma_rx_descriptor_slave_byteenable                        (mm_interconnect_0_sys_ethernet_dma_rx_descriptor_slave_byteenable),  //  output,   width = 32,                                                                 .byteenable
		.sys_ethernet_dma_rx_descriptor_slave_waitrequest                       (mm_interconnect_0_sys_ethernet_dma_rx_descriptor_slave_waitrequest), //   input,    width = 1,                                                                 .waitrequest
		.sys_ethernet_dma_tx_descriptor_slave_write                             (mm_interconnect_0_sys_ethernet_dma_tx_descriptor_slave_write),       //  output,    width = 1,                             sys_ethernet_dma_tx_descriptor_slave.write
		.sys_ethernet_dma_tx_descriptor_slave_writedata                         (mm_interconnect_0_sys_ethernet_dma_tx_descriptor_slave_writedata),   //  output,  width = 256,                                                                 .writedata
		.sys_ethernet_dma_tx_descriptor_slave_byteenable                        (mm_interconnect_0_sys_ethernet_dma_tx_descriptor_slave_byteenable),  //  output,   width = 32,                                                                 .byteenable
		.sys_ethernet_dma_tx_descriptor_slave_waitrequest                       (mm_interconnect_0_sys_ethernet_dma_tx_descriptor_slave_waitrequest), //   input,    width = 1,                                                                 .waitrequest
		.avl_adxcfg_0_rcfg_s0_address                                           (mm_interconnect_0_avl_adxcfg_0_rcfg_s0_address),                     //  output,   width = 10,                                             avl_adxcfg_0_rcfg_s0.address
		.avl_adxcfg_0_rcfg_s0_write                                             (mm_interconnect_0_avl_adxcfg_0_rcfg_s0_write),                       //  output,    width = 1,                                                                 .write
		.avl_adxcfg_0_rcfg_s0_read                                              (mm_interconnect_0_avl_adxcfg_0_rcfg_s0_read),                        //  output,    width = 1,                                                                 .read
		.avl_adxcfg_0_rcfg_s0_readdata                                          (mm_interconnect_0_avl_adxcfg_0_rcfg_s0_readdata),                    //   input,   width = 32,                                                                 .readdata
		.avl_adxcfg_0_rcfg_s0_writedata                                         (mm_interconnect_0_avl_adxcfg_0_rcfg_s0_writedata),                   //  output,   width = 32,                                                                 .writedata
		.avl_adxcfg_0_rcfg_s0_waitrequest                                       (mm_interconnect_0_avl_adxcfg_0_rcfg_s0_waitrequest),                 //   input,    width = 1,                                                                 .waitrequest
		.avl_adxcfg_1_rcfg_s0_address                                           (mm_interconnect_0_avl_adxcfg_1_rcfg_s0_address),                     //  output,   width = 10,                                             avl_adxcfg_1_rcfg_s0.address
		.avl_adxcfg_1_rcfg_s0_write                                             (mm_interconnect_0_avl_adxcfg_1_rcfg_s0_write),                       //  output,    width = 1,                                                                 .write
		.avl_adxcfg_1_rcfg_s0_read                                              (mm_interconnect_0_avl_adxcfg_1_rcfg_s0_read),                        //  output,    width = 1,                                                                 .read
		.avl_adxcfg_1_rcfg_s0_readdata                                          (mm_interconnect_0_avl_adxcfg_1_rcfg_s0_readdata),                    //   input,   width = 32,                                                                 .readdata
		.avl_adxcfg_1_rcfg_s0_writedata                                         (mm_interconnect_0_avl_adxcfg_1_rcfg_s0_writedata),                   //  output,   width = 32,                                                                 .writedata
		.avl_adxcfg_1_rcfg_s0_waitrequest                                       (mm_interconnect_0_avl_adxcfg_1_rcfg_s0_waitrequest),                 //   input,    width = 1,                                                                 .waitrequest
		.avl_adxcfg_2_rcfg_s0_address                                           (mm_interconnect_0_avl_adxcfg_2_rcfg_s0_address),                     //  output,   width = 10,                                             avl_adxcfg_2_rcfg_s0.address
		.avl_adxcfg_2_rcfg_s0_write                                             (mm_interconnect_0_avl_adxcfg_2_rcfg_s0_write),                       //  output,    width = 1,                                                                 .write
		.avl_adxcfg_2_rcfg_s0_read                                              (mm_interconnect_0_avl_adxcfg_2_rcfg_s0_read),                        //  output,    width = 1,                                                                 .read
		.avl_adxcfg_2_rcfg_s0_readdata                                          (mm_interconnect_0_avl_adxcfg_2_rcfg_s0_readdata),                    //   input,   width = 32,                                                                 .readdata
		.avl_adxcfg_2_rcfg_s0_writedata                                         (mm_interconnect_0_avl_adxcfg_2_rcfg_s0_writedata),                   //  output,   width = 32,                                                                 .writedata
		.avl_adxcfg_2_rcfg_s0_waitrequest                                       (mm_interconnect_0_avl_adxcfg_2_rcfg_s0_waitrequest),                 //   input,    width = 1,                                                                 .waitrequest
		.avl_adxcfg_3_rcfg_s0_address                                           (mm_interconnect_0_avl_adxcfg_3_rcfg_s0_address),                     //  output,   width = 10,                                             avl_adxcfg_3_rcfg_s0.address
		.avl_adxcfg_3_rcfg_s0_write                                             (mm_interconnect_0_avl_adxcfg_3_rcfg_s0_write),                       //  output,    width = 1,                                                                 .write
		.avl_adxcfg_3_rcfg_s0_read                                              (mm_interconnect_0_avl_adxcfg_3_rcfg_s0_read),                        //  output,    width = 1,                                                                 .read
		.avl_adxcfg_3_rcfg_s0_readdata                                          (mm_interconnect_0_avl_adxcfg_3_rcfg_s0_readdata),                    //   input,   width = 32,                                                                 .readdata
		.avl_adxcfg_3_rcfg_s0_writedata                                         (mm_interconnect_0_avl_adxcfg_3_rcfg_s0_writedata),                   //  output,   width = 32,                                                                 .writedata
		.avl_adxcfg_3_rcfg_s0_waitrequest                                       (mm_interconnect_0_avl_adxcfg_3_rcfg_s0_waitrequest),                 //   input,    width = 1,                                                                 .waitrequest
		.avl_adxcfg_0_rcfg_s1_address                                           (mm_interconnect_0_avl_adxcfg_0_rcfg_s1_address),                     //  output,   width = 10,                                             avl_adxcfg_0_rcfg_s1.address
		.avl_adxcfg_0_rcfg_s1_write                                             (mm_interconnect_0_avl_adxcfg_0_rcfg_s1_write),                       //  output,    width = 1,                                                                 .write
		.avl_adxcfg_0_rcfg_s1_read                                              (mm_interconnect_0_avl_adxcfg_0_rcfg_s1_read),                        //  output,    width = 1,                                                                 .read
		.avl_adxcfg_0_rcfg_s1_readdata                                          (mm_interconnect_0_avl_adxcfg_0_rcfg_s1_readdata),                    //   input,   width = 32,                                                                 .readdata
		.avl_adxcfg_0_rcfg_s1_writedata                                         (mm_interconnect_0_avl_adxcfg_0_rcfg_s1_writedata),                   //  output,   width = 32,                                                                 .writedata
		.avl_adxcfg_0_rcfg_s1_waitrequest                                       (mm_interconnect_0_avl_adxcfg_0_rcfg_s1_waitrequest),                 //   input,    width = 1,                                                                 .waitrequest
		.avl_adxcfg_1_rcfg_s1_address                                           (mm_interconnect_0_avl_adxcfg_1_rcfg_s1_address),                     //  output,   width = 10,                                             avl_adxcfg_1_rcfg_s1.address
		.avl_adxcfg_1_rcfg_s1_write                                             (mm_interconnect_0_avl_adxcfg_1_rcfg_s1_write),                       //  output,    width = 1,                                                                 .write
		.avl_adxcfg_1_rcfg_s1_read                                              (mm_interconnect_0_avl_adxcfg_1_rcfg_s1_read),                        //  output,    width = 1,                                                                 .read
		.avl_adxcfg_1_rcfg_s1_readdata                                          (mm_interconnect_0_avl_adxcfg_1_rcfg_s1_readdata),                    //   input,   width = 32,                                                                 .readdata
		.avl_adxcfg_1_rcfg_s1_writedata                                         (mm_interconnect_0_avl_adxcfg_1_rcfg_s1_writedata),                   //  output,   width = 32,                                                                 .writedata
		.avl_adxcfg_1_rcfg_s1_waitrequest                                       (mm_interconnect_0_avl_adxcfg_1_rcfg_s1_waitrequest),                 //   input,    width = 1,                                                                 .waitrequest
		.avl_adxcfg_2_rcfg_s1_address                                           (mm_interconnect_0_avl_adxcfg_2_rcfg_s1_address),                     //  output,   width = 10,                                             avl_adxcfg_2_rcfg_s1.address
		.avl_adxcfg_2_rcfg_s1_write                                             (mm_interconnect_0_avl_adxcfg_2_rcfg_s1_write),                       //  output,    width = 1,                                                                 .write
		.avl_adxcfg_2_rcfg_s1_read                                              (mm_interconnect_0_avl_adxcfg_2_rcfg_s1_read),                        //  output,    width = 1,                                                                 .read
		.avl_adxcfg_2_rcfg_s1_readdata                                          (mm_interconnect_0_avl_adxcfg_2_rcfg_s1_readdata),                    //   input,   width = 32,                                                                 .readdata
		.avl_adxcfg_2_rcfg_s1_writedata                                         (mm_interconnect_0_avl_adxcfg_2_rcfg_s1_writedata),                   //  output,   width = 32,                                                                 .writedata
		.avl_adxcfg_2_rcfg_s1_waitrequest                                       (mm_interconnect_0_avl_adxcfg_2_rcfg_s1_waitrequest),                 //   input,    width = 1,                                                                 .waitrequest
		.avl_adxcfg_3_rcfg_s1_address                                           (mm_interconnect_0_avl_adxcfg_3_rcfg_s1_address),                     //  output,   width = 10,                                             avl_adxcfg_3_rcfg_s1.address
		.avl_adxcfg_3_rcfg_s1_write                                             (mm_interconnect_0_avl_adxcfg_3_rcfg_s1_write),                       //  output,    width = 1,                                                                 .write
		.avl_adxcfg_3_rcfg_s1_read                                              (mm_interconnect_0_avl_adxcfg_3_rcfg_s1_read),                        //  output,    width = 1,                                                                 .read
		.avl_adxcfg_3_rcfg_s1_readdata                                          (mm_interconnect_0_avl_adxcfg_3_rcfg_s1_readdata),                    //   input,   width = 32,                                                                 .readdata
		.avl_adxcfg_3_rcfg_s1_writedata                                         (mm_interconnect_0_avl_adxcfg_3_rcfg_s1_writedata),                   //  output,   width = 32,                                                                 .writedata
		.avl_adxcfg_3_rcfg_s1_waitrequest                                       (mm_interconnect_0_avl_adxcfg_3_rcfg_s1_waitrequest),                 //   input,    width = 1,                                                                 .waitrequest
		.sys_ethernet_dma_rx_response_address                                   (mm_interconnect_0_sys_ethernet_dma_rx_response_address),             //  output,    width = 1,                                     sys_ethernet_dma_rx_response.address
		.sys_ethernet_dma_rx_response_read                                      (mm_interconnect_0_sys_ethernet_dma_rx_response_read),                //  output,    width = 1,                                                                 .read
		.sys_ethernet_dma_rx_response_readdata                                  (mm_interconnect_0_sys_ethernet_dma_rx_response_readdata),            //   input,   width = 32,                                                                 .readdata
		.sys_ethernet_dma_rx_response_byteenable                                (mm_interconnect_0_sys_ethernet_dma_rx_response_byteenable),          //  output,    width = 4,                                                                 .byteenable
		.sys_ethernet_dma_rx_response_waitrequest                               (mm_interconnect_0_sys_ethernet_dma_rx_response_waitrequest),         //   input,    width = 1,                                                                 .waitrequest
		.sys_int_mem_s1_address                                                 (mm_interconnect_0_sys_int_mem_s1_address),                           //  output,   width = 16,                                                   sys_int_mem_s1.address
		.sys_int_mem_s1_write                                                   (mm_interconnect_0_sys_int_mem_s1_write),                             //  output,    width = 1,                                                                 .write
		.sys_int_mem_s1_readdata                                                (mm_interconnect_0_sys_int_mem_s1_readdata),                          //   input,   width = 32,                                                                 .readdata
		.sys_int_mem_s1_writedata                                               (mm_interconnect_0_sys_int_mem_s1_writedata),                         //  output,   width = 32,                                                                 .writedata
		.sys_int_mem_s1_byteenable                                              (mm_interconnect_0_sys_int_mem_s1_byteenable),                        //  output,    width = 4,                                                                 .byteenable
		.sys_int_mem_s1_chipselect                                              (mm_interconnect_0_sys_int_mem_s1_chipselect),                        //  output,    width = 1,                                                                 .chipselect
		.sys_int_mem_s1_clken                                                   (mm_interconnect_0_sys_int_mem_s1_clken),                             //  output,    width = 1,                                                                 .clken
		.sys_timer_1_s1_address                                                 (mm_interconnect_0_sys_timer_1_s1_address),                           //  output,    width = 3,                                                   sys_timer_1_s1.address
		.sys_timer_1_s1_write                                                   (mm_interconnect_0_sys_timer_1_s1_write),                             //  output,    width = 1,                                                                 .write
		.sys_timer_1_s1_readdata                                                (mm_interconnect_0_sys_timer_1_s1_readdata),                          //   input,   width = 16,                                                                 .readdata
		.sys_timer_1_s1_writedata                                               (mm_interconnect_0_sys_timer_1_s1_writedata),                         //  output,   width = 16,                                                                 .writedata
		.sys_timer_1_s1_chipselect                                              (mm_interconnect_0_sys_timer_1_s1_chipselect),                        //  output,    width = 1,                                                                 .chipselect
		.sys_timer_2_s1_address                                                 (mm_interconnect_0_sys_timer_2_s1_address),                           //  output,    width = 3,                                                   sys_timer_2_s1.address
		.sys_timer_2_s1_write                                                   (mm_interconnect_0_sys_timer_2_s1_write),                             //  output,    width = 1,                                                                 .write
		.sys_timer_2_s1_readdata                                                (mm_interconnect_0_sys_timer_2_s1_readdata),                          //   input,   width = 16,                                                                 .readdata
		.sys_timer_2_s1_writedata                                               (mm_interconnect_0_sys_timer_2_s1_writedata),                         //  output,   width = 16,                                                                 .writedata
		.sys_timer_2_s1_chipselect                                              (mm_interconnect_0_sys_timer_2_s1_chipselect),                        //  output,    width = 1,                                                                 .chipselect
		.sys_gpio_bd_s1_address                                                 (mm_interconnect_0_sys_gpio_bd_s1_address),                           //  output,    width = 2,                                                   sys_gpio_bd_s1.address
		.sys_gpio_bd_s1_write                                                   (mm_interconnect_0_sys_gpio_bd_s1_write),                             //  output,    width = 1,                                                                 .write
		.sys_gpio_bd_s1_readdata                                                (mm_interconnect_0_sys_gpio_bd_s1_readdata),                          //   input,   width = 32,                                                                 .readdata
		.sys_gpio_bd_s1_writedata                                               (mm_interconnect_0_sys_gpio_bd_s1_writedata),                         //  output,   width = 32,                                                                 .writedata
		.sys_gpio_bd_s1_chipselect                                              (mm_interconnect_0_sys_gpio_bd_s1_chipselect),                        //  output,    width = 1,                                                                 .chipselect
		.sys_gpio_in_s1_address                                                 (mm_interconnect_0_sys_gpio_in_s1_address),                           //  output,    width = 2,                                                   sys_gpio_in_s1.address
		.sys_gpio_in_s1_write                                                   (mm_interconnect_0_sys_gpio_in_s1_write),                             //  output,    width = 1,                                                                 .write
		.sys_gpio_in_s1_readdata                                                (mm_interconnect_0_sys_gpio_in_s1_readdata),                          //   input,   width = 32,                                                                 .readdata
		.sys_gpio_in_s1_writedata                                               (mm_interconnect_0_sys_gpio_in_s1_writedata),                         //  output,   width = 32,                                                                 .writedata
		.sys_gpio_in_s1_chipselect                                              (mm_interconnect_0_sys_gpio_in_s1_chipselect),                        //  output,    width = 1,                                                                 .chipselect
		.sys_gpio_out_s1_address                                                (mm_interconnect_0_sys_gpio_out_s1_address),                          //  output,    width = 2,                                                  sys_gpio_out_s1.address
		.sys_gpio_out_s1_write                                                  (mm_interconnect_0_sys_gpio_out_s1_write),                            //  output,    width = 1,                                                                 .write
		.sys_gpio_out_s1_readdata                                               (mm_interconnect_0_sys_gpio_out_s1_readdata),                         //   input,   width = 32,                                                                 .readdata
		.sys_gpio_out_s1_writedata                                              (mm_interconnect_0_sys_gpio_out_s1_writedata),                        //  output,   width = 32,                                                                 .writedata
		.sys_gpio_out_s1_chipselect                                             (mm_interconnect_0_sys_gpio_out_s1_chipselect),                       //  output,    width = 1,                                                                 .chipselect
		.sys_spi_spi_control_port_address                                       (mm_interconnect_0_sys_spi_spi_control_port_address),                 //  output,    width = 3,                                         sys_spi_spi_control_port.address
		.sys_spi_spi_control_port_write                                         (mm_interconnect_0_sys_spi_spi_control_port_write),                   //  output,    width = 1,                                                                 .write
		.sys_spi_spi_control_port_read                                          (mm_interconnect_0_sys_spi_spi_control_port_read),                    //  output,    width = 1,                                                                 .read
		.sys_spi_spi_control_port_readdata                                      (mm_interconnect_0_sys_spi_spi_control_port_readdata),                //   input,   width = 16,                                                                 .readdata
		.sys_spi_spi_control_port_writedata                                     (mm_interconnect_0_sys_spi_spi_control_port_writedata),               //  output,   width = 16,                                                                 .writedata
		.sys_spi_spi_control_port_chipselect                                    (mm_interconnect_0_sys_spi_spi_control_port_chipselect),              //  output,    width = 1,                                                                 .chipselect
		.sys_flash_uas_address                                                  (mm_interconnect_0_sys_flash_uas_address),                            //  output,   width = 24,                                                    sys_flash_uas.address
		.sys_flash_uas_write                                                    (mm_interconnect_0_sys_flash_uas_write),                              //  output,    width = 1,                                                                 .write
		.sys_flash_uas_read                                                     (mm_interconnect_0_sys_flash_uas_read),                               //  output,    width = 1,                                                                 .read
		.sys_flash_uas_readdata                                                 (mm_interconnect_0_sys_flash_uas_readdata),                           //   input,   width = 32,                                                                 .readdata
		.sys_flash_uas_writedata                                                (mm_interconnect_0_sys_flash_uas_writedata),                          //  output,   width = 32,                                                                 .writedata
		.sys_flash_uas_burstcount                                               (mm_interconnect_0_sys_flash_uas_burstcount),                         //  output,    width = 3,                                                                 .burstcount
		.sys_flash_uas_byteenable                                               (mm_interconnect_0_sys_flash_uas_byteenable),                         //  output,    width = 4,                                                                 .byteenable
		.sys_flash_uas_readdatavalid                                            (mm_interconnect_0_sys_flash_uas_readdatavalid),                      //   input,    width = 1,                                                                 .readdatavalid
		.sys_flash_uas_waitrequest                                              (mm_interconnect_0_sys_flash_uas_waitrequest),                        //   input,    width = 1,                                                                 .waitrequest
		.sys_flash_uas_lock                                                     (mm_interconnect_0_sys_flash_uas_lock),                               //  output,    width = 1,                                                                 .lock
		.sys_flash_uas_debugaccess                                              (mm_interconnect_0_sys_flash_uas_debugaccess),                        //  output,    width = 1,                                                                 .debugaccess
		.axi_ad9680_dma_m_dest_axi_awid                                         (axi_ad9680_dma_m_dest_axi_awid),                                     //   input,    width = 1,                                        axi_ad9680_dma_m_dest_axi.awid
		.axi_ad9680_dma_m_dest_axi_awaddr                                       (axi_ad9680_dma_m_dest_axi_awaddr),                                   //   input,   width = 32,                                                                 .awaddr
		.axi_ad9680_dma_m_dest_axi_awlen                                        (axi_ad9680_dma_m_dest_axi_awlen),                                    //   input,    width = 4,                                                                 .awlen
		.axi_ad9680_dma_m_dest_axi_awsize                                       (axi_ad9680_dma_m_dest_axi_awsize),                                   //   input,    width = 3,                                                                 .awsize
		.axi_ad9680_dma_m_dest_axi_awburst                                      (axi_ad9680_dma_m_dest_axi_awburst),                                  //   input,    width = 2,                                                                 .awburst
		.axi_ad9680_dma_m_dest_axi_awlock                                       (axi_ad9680_dma_m_dest_axi_awlock),                                   //   input,    width = 2,                                                                 .awlock
		.axi_ad9680_dma_m_dest_axi_awcache                                      (axi_ad9680_dma_m_dest_axi_awcache),                                  //   input,    width = 4,                                                                 .awcache
		.axi_ad9680_dma_m_dest_axi_awprot                                       (axi_ad9680_dma_m_dest_axi_awprot),                                   //   input,    width = 3,                                                                 .awprot
		.axi_ad9680_dma_m_dest_axi_awvalid                                      (axi_ad9680_dma_m_dest_axi_awvalid),                                  //   input,    width = 1,                                                                 .awvalid
		.axi_ad9680_dma_m_dest_axi_awready                                      (axi_ad9680_dma_m_dest_axi_awready),                                  //  output,    width = 1,                                                                 .awready
		.axi_ad9680_dma_m_dest_axi_wid                                          (axi_ad9680_dma_m_dest_axi_wid),                                      //   input,    width = 1,                                                                 .wid
		.axi_ad9680_dma_m_dest_axi_wdata                                        (axi_ad9680_dma_m_dest_axi_wdata),                                    //   input,  width = 128,                                                                 .wdata
		.axi_ad9680_dma_m_dest_axi_wstrb                                        (axi_ad9680_dma_m_dest_axi_wstrb),                                    //   input,   width = 16,                                                                 .wstrb
		.axi_ad9680_dma_m_dest_axi_wlast                                        (axi_ad9680_dma_m_dest_axi_wlast),                                    //   input,    width = 1,                                                                 .wlast
		.axi_ad9680_dma_m_dest_axi_wvalid                                       (axi_ad9680_dma_m_dest_axi_wvalid),                                   //   input,    width = 1,                                                                 .wvalid
		.axi_ad9680_dma_m_dest_axi_wready                                       (axi_ad9680_dma_m_dest_axi_wready),                                   //  output,    width = 1,                                                                 .wready
		.axi_ad9680_dma_m_dest_axi_bid                                          (axi_ad9680_dma_m_dest_axi_bid),                                      //  output,    width = 1,                                                                 .bid
		.axi_ad9680_dma_m_dest_axi_bresp                                        (axi_ad9680_dma_m_dest_axi_bresp),                                    //  output,    width = 2,                                                                 .bresp
		.axi_ad9680_dma_m_dest_axi_bvalid                                       (axi_ad9680_dma_m_dest_axi_bvalid),                                   //  output,    width = 1,                                                                 .bvalid
		.axi_ad9680_dma_m_dest_axi_bready                                       (axi_ad9680_dma_m_dest_axi_bready),                                   //   input,    width = 1,                                                                 .bready
		.axi_ad9680_dma_m_dest_axi_arid                                         (axi_ad9680_dma_m_dest_axi_arid),                                     //   input,    width = 1,                                                                 .arid
		.axi_ad9680_dma_m_dest_axi_araddr                                       (axi_ad9680_dma_m_dest_axi_araddr),                                   //   input,   width = 32,                                                                 .araddr
		.axi_ad9680_dma_m_dest_axi_arlen                                        (axi_ad9680_dma_m_dest_axi_arlen),                                    //   input,    width = 4,                                                                 .arlen
		.axi_ad9680_dma_m_dest_axi_arsize                                       (axi_ad9680_dma_m_dest_axi_arsize),                                   //   input,    width = 3,                                                                 .arsize
		.axi_ad9680_dma_m_dest_axi_arburst                                      (axi_ad9680_dma_m_dest_axi_arburst),                                  //   input,    width = 2,                                                                 .arburst
		.axi_ad9680_dma_m_dest_axi_arlock                                       (axi_ad9680_dma_m_dest_axi_arlock),                                   //   input,    width = 2,                                                                 .arlock
		.axi_ad9680_dma_m_dest_axi_arcache                                      (axi_ad9680_dma_m_dest_axi_arcache),                                  //   input,    width = 4,                                                                 .arcache
		.axi_ad9680_dma_m_dest_axi_arprot                                       (axi_ad9680_dma_m_dest_axi_arprot),                                   //   input,    width = 3,                                                                 .arprot
		.axi_ad9680_dma_m_dest_axi_arvalid                                      (axi_ad9680_dma_m_dest_axi_arvalid),                                  //   input,    width = 1,                                                                 .arvalid
		.axi_ad9680_dma_m_dest_axi_arready                                      (axi_ad9680_dma_m_dest_axi_arready),                                  //  output,    width = 1,                                                                 .arready
		.axi_ad9680_dma_m_dest_axi_rid                                          (axi_ad9680_dma_m_dest_axi_rid),                                      //  output,    width = 1,                                                                 .rid
		.axi_ad9680_dma_m_dest_axi_rdata                                        (axi_ad9680_dma_m_dest_axi_rdata),                                    //  output,  width = 128,                                                                 .rdata
		.axi_ad9680_dma_m_dest_axi_rresp                                        (axi_ad9680_dma_m_dest_axi_rresp),                                    //  output,    width = 2,                                                                 .rresp
		.axi_ad9680_dma_m_dest_axi_rlast                                        (axi_ad9680_dma_m_dest_axi_rlast),                                    //  output,    width = 1,                                                                 .rlast
		.axi_ad9680_dma_m_dest_axi_rvalid                                       (axi_ad9680_dma_m_dest_axi_rvalid),                                   //  output,    width = 1,                                                                 .rvalid
		.axi_ad9680_dma_m_dest_axi_rready                                       (axi_ad9680_dma_m_dest_axi_rready),                                   //   input,    width = 1,                                                                 .rready
		.axi_ad9144_dma_m_src_axi_awid                                          (axi_ad9144_dma_m_src_axi_awid),                                      //   input,    width = 1,                                         axi_ad9144_dma_m_src_axi.awid
		.axi_ad9144_dma_m_src_axi_awaddr                                        (axi_ad9144_dma_m_src_axi_awaddr),                                    //   input,   width = 32,                                                                 .awaddr
		.axi_ad9144_dma_m_src_axi_awlen                                         (axi_ad9144_dma_m_src_axi_awlen),                                     //   input,    width = 4,                                                                 .awlen
		.axi_ad9144_dma_m_src_axi_awsize                                        (axi_ad9144_dma_m_src_axi_awsize),                                    //   input,    width = 3,                                                                 .awsize
		.axi_ad9144_dma_m_src_axi_awburst                                       (axi_ad9144_dma_m_src_axi_awburst),                                   //   input,    width = 2,                                                                 .awburst
		.axi_ad9144_dma_m_src_axi_awlock                                        (axi_ad9144_dma_m_src_axi_awlock),                                    //   input,    width = 2,                                                                 .awlock
		.axi_ad9144_dma_m_src_axi_awcache                                       (axi_ad9144_dma_m_src_axi_awcache),                                   //   input,    width = 4,                                                                 .awcache
		.axi_ad9144_dma_m_src_axi_awprot                                        (axi_ad9144_dma_m_src_axi_awprot),                                    //   input,    width = 3,                                                                 .awprot
		.axi_ad9144_dma_m_src_axi_awvalid                                       (axi_ad9144_dma_m_src_axi_awvalid),                                   //   input,    width = 1,                                                                 .awvalid
		.axi_ad9144_dma_m_src_axi_awready                                       (axi_ad9144_dma_m_src_axi_awready),                                   //  output,    width = 1,                                                                 .awready
		.axi_ad9144_dma_m_src_axi_wid                                           (axi_ad9144_dma_m_src_axi_wid),                                       //   input,    width = 1,                                                                 .wid
		.axi_ad9144_dma_m_src_axi_wdata                                         (axi_ad9144_dma_m_src_axi_wdata),                                     //   input,  width = 128,                                                                 .wdata
		.axi_ad9144_dma_m_src_axi_wstrb                                         (axi_ad9144_dma_m_src_axi_wstrb),                                     //   input,   width = 16,                                                                 .wstrb
		.axi_ad9144_dma_m_src_axi_wlast                                         (axi_ad9144_dma_m_src_axi_wlast),                                     //   input,    width = 1,                                                                 .wlast
		.axi_ad9144_dma_m_src_axi_wvalid                                        (axi_ad9144_dma_m_src_axi_wvalid),                                    //   input,    width = 1,                                                                 .wvalid
		.axi_ad9144_dma_m_src_axi_wready                                        (axi_ad9144_dma_m_src_axi_wready),                                    //  output,    width = 1,                                                                 .wready
		.axi_ad9144_dma_m_src_axi_bid                                           (axi_ad9144_dma_m_src_axi_bid),                                       //  output,    width = 1,                                                                 .bid
		.axi_ad9144_dma_m_src_axi_bresp                                         (axi_ad9144_dma_m_src_axi_bresp),                                     //  output,    width = 2,                                                                 .bresp
		.axi_ad9144_dma_m_src_axi_bvalid                                        (axi_ad9144_dma_m_src_axi_bvalid),                                    //  output,    width = 1,                                                                 .bvalid
		.axi_ad9144_dma_m_src_axi_bready                                        (axi_ad9144_dma_m_src_axi_bready),                                    //   input,    width = 1,                                                                 .bready
		.axi_ad9144_dma_m_src_axi_arid                                          (axi_ad9144_dma_m_src_axi_arid),                                      //   input,    width = 1,                                                                 .arid
		.axi_ad9144_dma_m_src_axi_araddr                                        (axi_ad9144_dma_m_src_axi_araddr),                                    //   input,   width = 32,                                                                 .araddr
		.axi_ad9144_dma_m_src_axi_arlen                                         (axi_ad9144_dma_m_src_axi_arlen),                                     //   input,    width = 4,                                                                 .arlen
		.axi_ad9144_dma_m_src_axi_arsize                                        (axi_ad9144_dma_m_src_axi_arsize),                                    //   input,    width = 3,                                                                 .arsize
		.axi_ad9144_dma_m_src_axi_arburst                                       (axi_ad9144_dma_m_src_axi_arburst),                                   //   input,    width = 2,                                                                 .arburst
		.axi_ad9144_dma_m_src_axi_arlock                                        (axi_ad9144_dma_m_src_axi_arlock),                                    //   input,    width = 2,                                                                 .arlock
		.axi_ad9144_dma_m_src_axi_arcache                                       (axi_ad9144_dma_m_src_axi_arcache),                                   //   input,    width = 4,                                                                 .arcache
		.axi_ad9144_dma_m_src_axi_arprot                                        (axi_ad9144_dma_m_src_axi_arprot),                                    //   input,    width = 3,                                                                 .arprot
		.axi_ad9144_dma_m_src_axi_arvalid                                       (axi_ad9144_dma_m_src_axi_arvalid),                                   //   input,    width = 1,                                                                 .arvalid
		.axi_ad9144_dma_m_src_axi_arready                                       (axi_ad9144_dma_m_src_axi_arready),                                   //  output,    width = 1,                                                                 .arready
		.axi_ad9144_dma_m_src_axi_rid                                           (axi_ad9144_dma_m_src_axi_rid),                                       //  output,    width = 1,                                                                 .rid
		.axi_ad9144_dma_m_src_axi_rdata                                         (axi_ad9144_dma_m_src_axi_rdata),                                     //  output,  width = 128,                                                                 .rdata
		.axi_ad9144_dma_m_src_axi_rresp                                         (axi_ad9144_dma_m_src_axi_rresp),                                     //  output,    width = 2,                                                                 .rresp
		.axi_ad9144_dma_m_src_axi_rlast                                         (axi_ad9144_dma_m_src_axi_rlast),                                     //  output,    width = 1,                                                                 .rlast
		.axi_ad9144_dma_m_src_axi_rvalid                                        (axi_ad9144_dma_m_src_axi_rvalid),                                    //  output,    width = 1,                                                                 .rvalid
		.axi_ad9144_dma_m_src_axi_rready                                        (axi_ad9144_dma_m_src_axi_rready),                                    //   input,    width = 1,                                                                 .rready
		.axi_ad9144_dma_s_axi_awaddr                                            (mm_interconnect_0_axi_ad9144_dma_s_axi_awaddr),                      //  output,   width = 12,                                             axi_ad9144_dma_s_axi.awaddr
		.axi_ad9144_dma_s_axi_awprot                                            (mm_interconnect_0_axi_ad9144_dma_s_axi_awprot),                      //  output,    width = 3,                                                                 .awprot
		.axi_ad9144_dma_s_axi_awvalid                                           (mm_interconnect_0_axi_ad9144_dma_s_axi_awvalid),                     //  output,    width = 1,                                                                 .awvalid
		.axi_ad9144_dma_s_axi_awready                                           (mm_interconnect_0_axi_ad9144_dma_s_axi_awready),                     //   input,    width = 1,                                                                 .awready
		.axi_ad9144_dma_s_axi_wdata                                             (mm_interconnect_0_axi_ad9144_dma_s_axi_wdata),                       //  output,   width = 32,                                                                 .wdata
		.axi_ad9144_dma_s_axi_wstrb                                             (mm_interconnect_0_axi_ad9144_dma_s_axi_wstrb),                       //  output,    width = 4,                                                                 .wstrb
		.axi_ad9144_dma_s_axi_wvalid                                            (mm_interconnect_0_axi_ad9144_dma_s_axi_wvalid),                      //  output,    width = 1,                                                                 .wvalid
		.axi_ad9144_dma_s_axi_wready                                            (mm_interconnect_0_axi_ad9144_dma_s_axi_wready),                      //   input,    width = 1,                                                                 .wready
		.axi_ad9144_dma_s_axi_bresp                                             (mm_interconnect_0_axi_ad9144_dma_s_axi_bresp),                       //   input,    width = 2,                                                                 .bresp
		.axi_ad9144_dma_s_axi_bvalid                                            (mm_interconnect_0_axi_ad9144_dma_s_axi_bvalid),                      //   input,    width = 1,                                                                 .bvalid
		.axi_ad9144_dma_s_axi_bready                                            (mm_interconnect_0_axi_ad9144_dma_s_axi_bready),                      //  output,    width = 1,                                                                 .bready
		.axi_ad9144_dma_s_axi_araddr                                            (mm_interconnect_0_axi_ad9144_dma_s_axi_araddr),                      //  output,   width = 12,                                                                 .araddr
		.axi_ad9144_dma_s_axi_arprot                                            (mm_interconnect_0_axi_ad9144_dma_s_axi_arprot),                      //  output,    width = 3,                                                                 .arprot
		.axi_ad9144_dma_s_axi_arvalid                                           (mm_interconnect_0_axi_ad9144_dma_s_axi_arvalid),                     //  output,    width = 1,                                                                 .arvalid
		.axi_ad9144_dma_s_axi_arready                                           (mm_interconnect_0_axi_ad9144_dma_s_axi_arready),                     //   input,    width = 1,                                                                 .arready
		.axi_ad9144_dma_s_axi_rdata                                             (mm_interconnect_0_axi_ad9144_dma_s_axi_rdata),                       //   input,   width = 32,                                                                 .rdata
		.axi_ad9144_dma_s_axi_rresp                                             (mm_interconnect_0_axi_ad9144_dma_s_axi_rresp),                       //   input,    width = 2,                                                                 .rresp
		.axi_ad9144_dma_s_axi_rvalid                                            (mm_interconnect_0_axi_ad9144_dma_s_axi_rvalid),                      //   input,    width = 1,                                                                 .rvalid
		.axi_ad9144_dma_s_axi_rready                                            (mm_interconnect_0_axi_ad9144_dma_s_axi_rready),                      //  output,    width = 1,                                                                 .rready
		.axi_ad9680_dma_s_axi_awaddr                                            (mm_interconnect_0_axi_ad9680_dma_s_axi_awaddr),                      //  output,   width = 12,                                             axi_ad9680_dma_s_axi.awaddr
		.axi_ad9680_dma_s_axi_awprot                                            (mm_interconnect_0_axi_ad9680_dma_s_axi_awprot),                      //  output,    width = 3,                                                                 .awprot
		.axi_ad9680_dma_s_axi_awvalid                                           (mm_interconnect_0_axi_ad9680_dma_s_axi_awvalid),                     //  output,    width = 1,                                                                 .awvalid
		.axi_ad9680_dma_s_axi_awready                                           (mm_interconnect_0_axi_ad9680_dma_s_axi_awready),                     //   input,    width = 1,                                                                 .awready
		.axi_ad9680_dma_s_axi_wdata                                             (mm_interconnect_0_axi_ad9680_dma_s_axi_wdata),                       //  output,   width = 32,                                                                 .wdata
		.axi_ad9680_dma_s_axi_wstrb                                             (mm_interconnect_0_axi_ad9680_dma_s_axi_wstrb),                       //  output,    width = 4,                                                                 .wstrb
		.axi_ad9680_dma_s_axi_wvalid                                            (mm_interconnect_0_axi_ad9680_dma_s_axi_wvalid),                      //  output,    width = 1,                                                                 .wvalid
		.axi_ad9680_dma_s_axi_wready                                            (mm_interconnect_0_axi_ad9680_dma_s_axi_wready),                      //   input,    width = 1,                                                                 .wready
		.axi_ad9680_dma_s_axi_bresp                                             (mm_interconnect_0_axi_ad9680_dma_s_axi_bresp),                       //   input,    width = 2,                                                                 .bresp
		.axi_ad9680_dma_s_axi_bvalid                                            (mm_interconnect_0_axi_ad9680_dma_s_axi_bvalid),                      //   input,    width = 1,                                                                 .bvalid
		.axi_ad9680_dma_s_axi_bready                                            (mm_interconnect_0_axi_ad9680_dma_s_axi_bready),                      //  output,    width = 1,                                                                 .bready
		.axi_ad9680_dma_s_axi_araddr                                            (mm_interconnect_0_axi_ad9680_dma_s_axi_araddr),                      //  output,   width = 12,                                                                 .araddr
		.axi_ad9680_dma_s_axi_arprot                                            (mm_interconnect_0_axi_ad9680_dma_s_axi_arprot),                      //  output,    width = 3,                                                                 .arprot
		.axi_ad9680_dma_s_axi_arvalid                                           (mm_interconnect_0_axi_ad9680_dma_s_axi_arvalid),                     //  output,    width = 1,                                                                 .arvalid
		.axi_ad9680_dma_s_axi_arready                                           (mm_interconnect_0_axi_ad9680_dma_s_axi_arready),                     //   input,    width = 1,                                                                 .arready
		.axi_ad9680_dma_s_axi_rdata                                             (mm_interconnect_0_axi_ad9680_dma_s_axi_rdata),                       //   input,   width = 32,                                                                 .rdata
		.axi_ad9680_dma_s_axi_rresp                                             (mm_interconnect_0_axi_ad9680_dma_s_axi_rresp),                       //   input,    width = 2,                                                                 .rresp
		.axi_ad9680_dma_s_axi_rvalid                                            (mm_interconnect_0_axi_ad9680_dma_s_axi_rvalid),                      //   input,    width = 1,                                                                 .rvalid
		.axi_ad9680_dma_s_axi_rready                                            (mm_interconnect_0_axi_ad9680_dma_s_axi_rready),                      //  output,    width = 1,                                                                 .rready
		.sys_cpu_reset_reset_bridge_in_reset_reset                              (rst_controller_004_reset_out_reset),                                 //   input,    width = 1,                              sys_cpu_reset_reset_bridge_in_reset.reset
		.axi_ad9680_dma_m_dest_axi_reset_reset_bridge_in_reset_reset            (rst_controller_002_reset_out_reset),                                 //   input,    width = 1,            axi_ad9680_dma_m_dest_axi_reset_reset_bridge_in_reset.reset
		.axi_ad9680_dma_s_axi_reset_reset_bridge_in_reset_reset                 (rst_controller_reset_out_reset),                                     //   input,    width = 1,                 axi_ad9680_dma_s_axi_reset_reset_bridge_in_reset.reset
		.sys_ddr3_cntrl_ctrl_amm_0_translator_reset_reset_bridge_in_reset_reset (rst_controller_006_reset_out_reset),                                 //   input,    width = 1, sys_ddr3_cntrl_ctrl_amm_0_translator_reset_reset_bridge_in_reset.reset
		.sys_clk_clk_clk                                                        (sys_clk_clk_clk),                                                    //   input,    width = 1,                                                      sys_clk_clk.clk
		.sys_ddr3_cntrl_emif_usr_clk_clk                                        (sys_ddr3_cntrl_emif_usr_clk_clk)                                     //   input,    width = 1,                                      sys_ddr3_cntrl_emif_usr_clk.clk
	);

	system_bd_altera_mm_interconnect_181_bnruudi mm_interconnect_1 (
		.sys_cpu_tightly_coupled_data_master_0_address    (sys_cpu_tightly_coupled_data_master_0_address),    //   input,  width = 29,    sys_cpu_tightly_coupled_data_master_0.address
		.sys_cpu_tightly_coupled_data_master_0_byteenable (sys_cpu_tightly_coupled_data_master_0_byteenable), //   input,   width = 4,                                         .byteenable
		.sys_cpu_tightly_coupled_data_master_0_read       (sys_cpu_tightly_coupled_data_master_0_read),       //   input,   width = 1,                                         .read
		.sys_cpu_tightly_coupled_data_master_0_readdata   (sys_cpu_tightly_coupled_data_master_0_readdata),   //  output,  width = 32,                                         .readdata
		.sys_cpu_tightly_coupled_data_master_0_write      (sys_cpu_tightly_coupled_data_master_0_write),      //   input,   width = 1,                                         .write
		.sys_cpu_tightly_coupled_data_master_0_writedata  (sys_cpu_tightly_coupled_data_master_0_writedata),  //   input,  width = 32,                                         .writedata
		.sys_tlb_mem_s1_address                           (mm_interconnect_1_sys_tlb_mem_s1_address),         //  output,  width = 16,                           sys_tlb_mem_s1.address
		.sys_tlb_mem_s1_write                             (mm_interconnect_1_sys_tlb_mem_s1_write),           //  output,   width = 1,                                         .write
		.sys_tlb_mem_s1_readdata                          (mm_interconnect_1_sys_tlb_mem_s1_readdata),        //   input,  width = 32,                                         .readdata
		.sys_tlb_mem_s1_writedata                         (mm_interconnect_1_sys_tlb_mem_s1_writedata),       //  output,  width = 32,                                         .writedata
		.sys_tlb_mem_s1_byteenable                        (mm_interconnect_1_sys_tlb_mem_s1_byteenable),      //  output,   width = 4,                                         .byteenable
		.sys_tlb_mem_s1_chipselect                        (mm_interconnect_1_sys_tlb_mem_s1_chipselect),      //  output,   width = 1,                                         .chipselect
		.sys_tlb_mem_s1_clken                             (mm_interconnect_1_sys_tlb_mem_s1_clken),           //  output,   width = 1,                                         .clken
		.sys_cpu_reset_reset_bridge_in_reset_reset        (rst_controller_004_reset_out_reset),               //   input,   width = 1,      sys_cpu_reset_reset_bridge_in_reset.reset
		.sys_tlb_mem_reset1_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                   //   input,   width = 1, sys_tlb_mem_reset1_reset_bridge_in_reset.reset
		.sys_clk_clk_clk                                  (sys_clk_clk_clk)                                   //   input,   width = 1,                              sys_clk_clk.clk
	);

	system_bd_altera_mm_interconnect_181_nxa5mji mm_interconnect_2 (
		.sys_cpu_tightly_coupled_instruction_master_0_address  (sys_cpu_tightly_coupled_instruction_master_0_address),  //   input,  width = 29, sys_cpu_tightly_coupled_instruction_master_0.address
		.sys_cpu_tightly_coupled_instruction_master_0_read     (sys_cpu_tightly_coupled_instruction_master_0_read),     //   input,   width = 1,                                             .read
		.sys_cpu_tightly_coupled_instruction_master_0_readdata (sys_cpu_tightly_coupled_instruction_master_0_readdata), //  output,  width = 32,                                             .readdata
		.sys_tlb_mem_s2_address                                (mm_interconnect_2_sys_tlb_mem_s2_address),              //  output,  width = 16,                               sys_tlb_mem_s2.address
		.sys_tlb_mem_s2_write                                  (mm_interconnect_2_sys_tlb_mem_s2_write),                //  output,   width = 1,                                             .write
		.sys_tlb_mem_s2_readdata                               (mm_interconnect_2_sys_tlb_mem_s2_readdata),             //   input,  width = 32,                                             .readdata
		.sys_tlb_mem_s2_writedata                              (mm_interconnect_2_sys_tlb_mem_s2_writedata),            //  output,  width = 32,                                             .writedata
		.sys_tlb_mem_s2_byteenable                             (mm_interconnect_2_sys_tlb_mem_s2_byteenable),           //  output,   width = 4,                                             .byteenable
		.sys_tlb_mem_s2_chipselect                             (mm_interconnect_2_sys_tlb_mem_s2_chipselect),           //  output,   width = 1,                                             .chipselect
		.sys_tlb_mem_s2_clken                                  (mm_interconnect_2_sys_tlb_mem_s2_clken),                //  output,   width = 1,                                             .clken
		.sys_cpu_reset_reset_bridge_in_reset_reset             (rst_controller_004_reset_out_reset),                    //   input,   width = 1,          sys_cpu_reset_reset_bridge_in_reset.reset
		.sys_tlb_mem_reset2_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                        //   input,   width = 1,     sys_tlb_mem_reset2_reset_bridge_in_reset.reset
		.sys_clk_clk_clk                                       (sys_clk_clk_clk)                                        //   input,   width = 1,                                  sys_clk_clk.clk
	);

	system_bd_altera_irq_mapper_181_zfhtbja irq_mapper (
		.clk           (sys_clk_clk_clk),                    //   input,   width = 1,       clk.clk
		.reset         (rst_controller_004_reset_out_reset), //   input,   width = 1, clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           //   input,   width = 1, receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           //   input,   width = 1, receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           //   input,   width = 1, receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           //   input,   width = 1, receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           //   input,   width = 1, receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           //   input,   width = 1, receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           //   input,   width = 1, receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),           //   input,   width = 1, receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),           //   input,   width = 1, receiver8.irq
		.receiver9_irq (irq_mapper_receiver9_irq),           //   input,   width = 1, receiver9.irq
		.sender_irq    (sys_cpu_irq_irq)                     //  output,  width = 32,    sender.irq
	);

	system_bd_altera_avalon_st_adapter_181_ffpp76a #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (6),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (sys_clk_clk_clk),                       //   input,   width = 1, in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),        //   input,   width = 1, in_rst_0.reset
		.out_0_data          (avalon_st_adapter_out_0_data),          //  output,  width = 64,    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //  output,   width = 1,         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //   input,   width = 1,         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //  output,   width = 1,         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //  output,   width = 1,         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //  output,   width = 3,         .empty
		.out_0_error         (avalon_st_adapter_out_0_error),         //  output,   width = 6,         .error
		.in_0_data           (sys_ethernet_receive_data),             //   input,  width = 32,     in_0.data
		.in_0_valid          (sys_ethernet_receive_valid),            //   input,   width = 1,         .valid
		.in_0_ready          (sys_ethernet_receive_ready),            //  output,   width = 1,         .ready
		.in_0_startofpacket  (sys_ethernet_receive_startofpacket),    //   input,   width = 1,         .startofpacket
		.in_0_endofpacket    (sys_ethernet_receive_endofpacket),      //   input,   width = 1,         .endofpacket
		.in_0_empty          (sys_ethernet_receive_empty),            //   input,   width = 2,         .empty
		.in_0_error          (sys_ethernet_receive_error)             //   input,   width = 6,         .error
	);

	system_bd_altera_avalon_st_adapter_181_r34pkoa #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (0),
		.inErrorWidth    (1),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (sys_clk_clk_clk),                             //   input,   width = 1, in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),              //   input,   width = 1, in_rst_0.reset
		.in_0_data           (sys_ethernet_dma_tx_st_source_data),          //   input,  width = 64,     in_0.data
		.in_0_valid          (sys_ethernet_dma_tx_st_source_valid),         //   input,   width = 1,         .valid
		.in_0_ready          (sys_ethernet_dma_tx_st_source_ready),         //  output,   width = 1,         .ready
		.in_0_startofpacket  (sys_ethernet_dma_tx_st_source_startofpacket), //   input,   width = 1,         .startofpacket
		.in_0_endofpacket    (sys_ethernet_dma_tx_st_source_endofpacket),   //   input,   width = 1,         .endofpacket
		.in_0_empty          (sys_ethernet_dma_tx_st_source_empty),         //   input,   width = 3,         .empty
		.in_0_error          (sys_ethernet_dma_tx_st_source_error),         //   input,   width = 1,         .error
		.out_0_data          (avalon_st_adapter_001_out_0_data),            //  output,  width = 32,    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),           //  output,   width = 1,         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),           //   input,   width = 1,         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket),   //  output,   width = 1,         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),     //  output,   width = 1,         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty),           //  output,   width = 2,         .empty
		.out_0_error         (avalon_st_adapter_001_out_0_error)            //  output,   width = 1,         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~sys_clk_clk_reset_reset),           //   input,  width = 1, reset_in0.reset
		.clk            (sys_clk_clk_clk),                    //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~sys_clk_clk_reset_reset),           //   input,  width = 1, reset_in0.reset
		.reset_in1      (~sys_dma_clk_clk_reset_reset),       //   input,  width = 1, reset_in1.reset
		.clk            (ad9680_jesd204_link_clk_clk),        //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~sys_dma_clk_clk_reset_reset),       //   input,  width = 1, reset_in0.reset
		.clk            (sys_ddr3_cntrl_emif_usr_clk_clk),    //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (ad9144_jesd204_link_reset_reset),    //   input,  width = 1, reset_in0.reset
		.clk            (ad9144_jesd204_link_clk_clk),        //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~sys_clk_clk_reset_reset),               //   input,  width = 1, reset_in0.reset
		.reset_in1      (sys_cpu_debug_reset_request_reset),      //   input,  width = 1, reset_in1.reset
		.clk            (sys_clk_clk_clk),                        //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_004_reset_out_reset_req), //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated),                       
		.reset_req_in1  (1'b0),                                   // (terminated),                       
		.reset_in2      (1'b0),                                   // (terminated),                       
		.reset_req_in2  (1'b0),                                   // (terminated),                       
		.reset_in3      (1'b0),                                   // (terminated),                       
		.reset_req_in3  (1'b0),                                   // (terminated),                       
		.reset_in4      (1'b0),                                   // (terminated),                       
		.reset_req_in4  (1'b0),                                   // (terminated),                       
		.reset_in5      (1'b0),                                   // (terminated),                       
		.reset_req_in5  (1'b0),                                   // (terminated),                       
		.reset_in6      (1'b0),                                   // (terminated),                       
		.reset_req_in6  (1'b0),                                   // (terminated),                       
		.reset_in7      (1'b0),                                   // (terminated),                       
		.reset_req_in7  (1'b0),                                   // (terminated),                       
		.reset_in8      (1'b0),                                   // (terminated),                       
		.reset_req_in8  (1'b0),                                   // (terminated),                       
		.reset_in9      (1'b0),                                   // (terminated),                       
		.reset_req_in9  (1'b0),                                   // (terminated),                       
		.reset_in10     (1'b0),                                   // (terminated),                       
		.reset_req_in10 (1'b0),                                   // (terminated),                       
		.reset_in11     (1'b0),                                   // (terminated),                       
		.reset_req_in11 (1'b0),                                   // (terminated),                       
		.reset_in12     (1'b0),                                   // (terminated),                       
		.reset_req_in12 (1'b0),                                   // (terminated),                       
		.reset_in13     (1'b0),                                   // (terminated),                       
		.reset_req_in13 (1'b0),                                   // (terminated),                       
		.reset_in14     (1'b0),                                   // (terminated),                       
		.reset_req_in14 (1'b0),                                   // (terminated),                       
		.reset_in15     (1'b0),                                   // (terminated),                       
		.reset_req_in15 (1'b0)                                    // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~sys_clk_clk_reset_reset),           //   input,  width = 1, reset_in0.reset
		.clk            (sys_clk_clk_clk),                    //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~sys_ddr3_cntrl_emif_usr_reset_n_reset), //   input,  width = 1, reset_in0.reset
		.clk            (sys_ddr3_cntrl_emif_usr_clk_clk),        //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (),                                       // (terminated),                       
		.reset_req_in0  (1'b0),                                   // (terminated),                       
		.reset_in1      (1'b0),                                   // (terminated),                       
		.reset_req_in1  (1'b0),                                   // (terminated),                       
		.reset_in2      (1'b0),                                   // (terminated),                       
		.reset_req_in2  (1'b0),                                   // (terminated),                       
		.reset_in3      (1'b0),                                   // (terminated),                       
		.reset_req_in3  (1'b0),                                   // (terminated),                       
		.reset_in4      (1'b0),                                   // (terminated),                       
		.reset_req_in4  (1'b0),                                   // (terminated),                       
		.reset_in5      (1'b0),                                   // (terminated),                       
		.reset_req_in5  (1'b0),                                   // (terminated),                       
		.reset_in6      (1'b0),                                   // (terminated),                       
		.reset_req_in6  (1'b0),                                   // (terminated),                       
		.reset_in7      (1'b0),                                   // (terminated),                       
		.reset_req_in7  (1'b0),                                   // (terminated),                       
		.reset_in8      (1'b0),                                   // (terminated),                       
		.reset_req_in8  (1'b0),                                   // (terminated),                       
		.reset_in9      (1'b0),                                   // (terminated),                       
		.reset_req_in9  (1'b0),                                   // (terminated),                       
		.reset_in10     (1'b0),                                   // (terminated),                       
		.reset_req_in10 (1'b0),                                   // (terminated),                       
		.reset_in11     (1'b0),                                   // (terminated),                       
		.reset_req_in11 (1'b0),                                   // (terminated),                       
		.reset_in12     (1'b0),                                   // (terminated),                       
		.reset_req_in12 (1'b0),                                   // (terminated),                       
		.reset_in13     (1'b0),                                   // (terminated),                       
		.reset_req_in13 (1'b0),                                   // (terminated),                       
		.reset_in14     (1'b0),                                   // (terminated),                       
		.reset_req_in14 (1'b0),                                   // (terminated),                       
		.reset_in15     (1'b0),                                   // (terminated),                       
		.reset_req_in15 (1'b0)                                    // (terminated),                       
	);

endmodule
